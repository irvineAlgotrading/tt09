magic
tech sky130B
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -91 6704 13433 7006
rect 1713 4527 13433 6704
rect 1713 4020 3576 4527
rect -91 3718 3576 4020
rect 18928 852 19259 2337
<< pwell >>
rect 13008 2834 19221 3039
rect 13008 1452 13657 2834
rect 15119 2776 19221 2834
rect 18988 2412 19221 2776
rect 10593 1366 13657 1452
rect 10593 1302 10679 1366
rect 10593 354 10679 478
rect 10593 320 15123 354
rect 19026 320 19180 790
rect 10593 64 19180 320
rect 18846 38 19180 64
<< mvpsubdiff >>
rect 13034 2979 13058 3013
rect 13092 2979 13127 3013
rect 13161 2979 13196 3013
rect 13230 2979 13265 3013
rect 13299 2979 13334 3013
rect 13368 2979 13403 3013
rect 13437 2979 13472 3013
rect 13506 2979 13541 3013
rect 13575 2979 13610 3013
rect 13644 2979 13679 3013
rect 13713 2979 13748 3013
rect 13782 2979 13817 3013
rect 13851 2979 13886 3013
rect 13920 2979 13955 3013
rect 13989 2979 14024 3013
rect 14058 2979 14093 3013
rect 14127 2979 14162 3013
rect 14196 2979 14231 3013
rect 14265 2979 14299 3013
rect 14333 2979 14367 3013
rect 14401 2979 14435 3013
rect 14469 2979 14503 3013
rect 14537 2979 14571 3013
rect 14605 2979 14639 3013
rect 14673 2979 14707 3013
rect 14741 2979 14775 3013
rect 14809 2979 14843 3013
rect 14877 2979 14911 3013
rect 14945 2979 14979 3013
rect 15013 2979 15047 3013
rect 15081 2979 15115 3013
rect 15149 2979 15183 3013
rect 15217 2979 15251 3013
rect 15285 2979 15319 3013
rect 15353 2979 15387 3013
rect 15421 2979 15455 3013
rect 15489 2979 15523 3013
rect 15557 2979 15591 3013
rect 15625 2979 15659 3013
rect 15693 2979 15727 3013
rect 15761 2979 15795 3013
rect 15829 2979 15863 3013
rect 15897 2979 15931 3013
rect 15965 2979 15999 3013
rect 16033 2979 16067 3013
rect 16101 2979 16135 3013
rect 16169 2979 16203 3013
rect 16237 2979 16271 3013
rect 16305 2979 16339 3013
rect 16373 2979 16407 3013
rect 16441 2979 16475 3013
rect 16509 2979 16543 3013
rect 16577 2979 16611 3013
rect 16645 2979 16679 3013
rect 16713 2979 16747 3013
rect 16781 2979 16815 3013
rect 16849 2979 16883 3013
rect 16917 2979 16951 3013
rect 16985 2979 17019 3013
rect 17053 2979 17087 3013
rect 17121 2979 17155 3013
rect 17189 2979 17223 3013
rect 17257 2979 17291 3013
rect 17325 2979 17359 3013
rect 17393 2979 17427 3013
rect 17461 2979 17495 3013
rect 17529 2979 17563 3013
rect 17597 2979 17631 3013
rect 17665 2979 17699 3013
rect 17733 2979 17767 3013
rect 17801 2979 17835 3013
rect 17869 2979 17903 3013
rect 17937 2979 17971 3013
rect 18005 2979 18039 3013
rect 19025 2979 19195 3013
rect 13034 2945 18067 2979
rect 19025 2945 19093 2979
rect 19127 2945 19195 2979
rect 13034 2911 15169 2945
rect 15203 2911 15238 2945
rect 15272 2911 15307 2945
rect 15341 2911 15376 2945
rect 15410 2911 15445 2945
rect 15479 2911 15514 2945
rect 15548 2911 15583 2945
rect 15617 2911 15652 2945
rect 15686 2911 15721 2945
rect 15755 2911 15790 2945
rect 15824 2911 15859 2945
rect 15893 2911 15928 2945
rect 15962 2911 15997 2945
rect 16031 2911 16066 2945
rect 16100 2911 16135 2945
rect 16169 2911 16204 2945
rect 16238 2911 16273 2945
rect 16307 2911 16342 2945
rect 16376 2911 16411 2945
rect 16445 2911 16480 2945
rect 16514 2911 16549 2945
rect 16583 2911 16618 2945
rect 16652 2911 16687 2945
rect 16721 2911 16756 2945
rect 16790 2911 16825 2945
rect 16859 2911 16894 2945
rect 16928 2911 16963 2945
rect 16997 2911 17032 2945
rect 17066 2911 17101 2945
rect 17135 2911 17170 2945
rect 17204 2911 17239 2945
rect 17273 2911 17308 2945
rect 17342 2911 17377 2945
rect 17411 2911 17446 2945
rect 17480 2911 17515 2945
rect 17549 2911 17584 2945
rect 17618 2911 17653 2945
rect 17687 2911 17722 2945
rect 17756 2911 17791 2945
rect 17825 2911 17860 2945
rect 17894 2911 17929 2945
rect 17963 2911 17998 2945
rect 18032 2911 18067 2945
rect 13034 2877 13058 2911
rect 13092 2877 13127 2911
rect 13161 2877 13196 2911
rect 13230 2877 13265 2911
rect 13299 2877 13334 2911
rect 13368 2877 13403 2911
rect 13437 2877 13472 2911
rect 13506 2877 13541 2911
rect 13575 2877 13610 2911
rect 13644 2877 13679 2911
rect 13713 2877 13748 2911
rect 13782 2877 13817 2911
rect 13851 2877 13886 2911
rect 13920 2877 13954 2911
rect 13988 2877 14022 2911
rect 14056 2877 14090 2911
rect 14124 2877 14158 2911
rect 14192 2877 14226 2911
rect 14260 2877 14294 2911
rect 14328 2877 14362 2911
rect 14396 2877 14430 2911
rect 14464 2877 14498 2911
rect 14532 2877 14566 2911
rect 14600 2877 14634 2911
rect 14668 2877 14702 2911
rect 14736 2877 14770 2911
rect 14804 2877 14838 2911
rect 14872 2877 14906 2911
rect 14940 2877 14974 2911
rect 15008 2877 15042 2911
rect 15076 2877 18067 2911
rect 13034 2860 15169 2877
rect 13034 2809 13631 2860
rect 13034 2775 13058 2809
rect 13092 2775 13126 2809
rect 13160 2775 13194 2809
rect 13228 2775 13262 2809
rect 13296 2775 13330 2809
rect 13364 2775 13398 2809
rect 13432 2775 13466 2809
rect 13500 2775 13631 2809
rect 15145 2843 15169 2860
rect 15203 2843 15238 2877
rect 15272 2843 15307 2877
rect 15341 2843 15376 2877
rect 15410 2843 15445 2877
rect 15479 2843 15514 2877
rect 15548 2843 15583 2877
rect 15617 2843 15652 2877
rect 15686 2843 15721 2877
rect 15755 2843 15790 2877
rect 15824 2843 15859 2877
rect 15893 2843 15928 2877
rect 15962 2843 15997 2877
rect 16031 2843 16066 2877
rect 16100 2843 16135 2877
rect 16169 2843 16204 2877
rect 16238 2843 16273 2877
rect 16307 2843 16342 2877
rect 16376 2843 16411 2877
rect 16445 2843 16480 2877
rect 16514 2843 16549 2877
rect 16583 2843 16618 2877
rect 16652 2843 16687 2877
rect 16721 2843 16756 2877
rect 16790 2843 16825 2877
rect 16859 2843 16894 2877
rect 16928 2843 16963 2877
rect 16997 2843 17032 2877
rect 17066 2843 17101 2877
rect 17135 2843 17170 2877
rect 17204 2843 17239 2877
rect 17273 2843 17308 2877
rect 17342 2843 17377 2877
rect 17411 2843 17446 2877
rect 17480 2843 17515 2877
rect 17549 2843 17584 2877
rect 17618 2843 17653 2877
rect 17687 2843 17722 2877
rect 17756 2843 17791 2877
rect 17825 2843 17860 2877
rect 17894 2843 17929 2877
rect 17963 2843 17998 2877
rect 18032 2843 18067 2877
rect 19053 2910 19195 2945
rect 19053 2876 19093 2910
rect 19127 2876 19195 2910
rect 19053 2843 19195 2876
rect 15145 2841 19195 2843
rect 15145 2807 19093 2841
rect 19127 2807 19195 2841
rect 15145 2802 19195 2807
rect 13034 2739 13631 2775
rect 13034 2705 13058 2739
rect 13092 2705 13126 2739
rect 13160 2705 13194 2739
rect 13228 2705 13262 2739
rect 13296 2705 13330 2739
rect 13364 2705 13398 2739
rect 13432 2705 13466 2739
rect 13500 2705 13631 2739
rect 13034 2669 13631 2705
rect 13034 2635 13058 2669
rect 13092 2635 13126 2669
rect 13160 2635 13194 2669
rect 13228 2635 13262 2669
rect 13296 2635 13330 2669
rect 13364 2635 13398 2669
rect 13432 2635 13466 2669
rect 13500 2635 13631 2669
rect 13034 2599 13631 2635
rect 13034 2565 13058 2599
rect 13092 2565 13126 2599
rect 13160 2565 13194 2599
rect 13228 2565 13262 2599
rect 13296 2565 13330 2599
rect 13364 2565 13398 2599
rect 13432 2565 13466 2599
rect 13500 2565 13631 2599
rect 13034 2529 13631 2565
rect 13034 2495 13058 2529
rect 13092 2495 13126 2529
rect 13160 2495 13194 2529
rect 13228 2495 13262 2529
rect 13296 2495 13330 2529
rect 13364 2495 13398 2529
rect 13432 2495 13466 2529
rect 13500 2495 13631 2529
rect 13034 2460 13631 2495
rect 13034 2426 13058 2460
rect 13092 2426 13126 2460
rect 13160 2426 13194 2460
rect 13228 2426 13262 2460
rect 13296 2426 13330 2460
rect 13364 2426 13398 2460
rect 13432 2426 13466 2460
rect 13500 2426 13631 2460
rect 19014 2772 19195 2802
rect 19014 2738 19093 2772
rect 19127 2738 19195 2772
rect 19014 2703 19195 2738
rect 19014 2669 19093 2703
rect 19127 2669 19195 2703
rect 19014 2634 19195 2669
rect 19014 2600 19093 2634
rect 19127 2600 19195 2634
rect 19014 2565 19195 2600
rect 19014 2531 19093 2565
rect 19127 2531 19195 2565
rect 19014 2496 19195 2531
rect 19014 2462 19093 2496
rect 19127 2462 19195 2496
rect 19014 2438 19195 2462
rect 13034 2391 13631 2426
rect 13034 2357 13058 2391
rect 13092 2357 13126 2391
rect 13160 2357 13194 2391
rect 13228 2357 13262 2391
rect 13296 2357 13330 2391
rect 13364 2357 13398 2391
rect 13432 2357 13466 2391
rect 13500 2357 13631 2391
rect 13034 2322 13631 2357
rect 13034 2288 13058 2322
rect 13092 2288 13126 2322
rect 13160 2288 13194 2322
rect 13228 2288 13262 2322
rect 13296 2288 13330 2322
rect 13364 2288 13398 2322
rect 13432 2288 13466 2322
rect 13500 2288 13631 2322
rect 13034 2253 13631 2288
rect 13034 2219 13058 2253
rect 13092 2219 13126 2253
rect 13160 2219 13194 2253
rect 13228 2219 13262 2253
rect 13296 2219 13330 2253
rect 13364 2219 13398 2253
rect 13432 2219 13466 2253
rect 13500 2219 13631 2253
rect 13034 2184 13631 2219
rect 13034 2150 13058 2184
rect 13092 2150 13126 2184
rect 13160 2150 13194 2184
rect 13228 2150 13262 2184
rect 13296 2150 13330 2184
rect 13364 2150 13398 2184
rect 13432 2150 13466 2184
rect 13500 2150 13631 2184
rect 13034 2115 13631 2150
rect 13034 2081 13058 2115
rect 13092 2081 13126 2115
rect 13160 2081 13194 2115
rect 13228 2081 13262 2115
rect 13296 2081 13330 2115
rect 13364 2081 13398 2115
rect 13432 2081 13466 2115
rect 13500 2081 13631 2115
rect 13034 2046 13631 2081
rect 13034 2012 13058 2046
rect 13092 2012 13126 2046
rect 13160 2012 13194 2046
rect 13228 2012 13262 2046
rect 13296 2012 13330 2046
rect 13364 2012 13398 2046
rect 13432 2012 13466 2046
rect 13500 2012 13631 2046
rect 13034 1977 13631 2012
rect 13034 1943 13058 1977
rect 13092 1943 13126 1977
rect 13160 1943 13194 1977
rect 13228 1943 13262 1977
rect 13296 1943 13330 1977
rect 13364 1943 13398 1977
rect 13432 1943 13466 1977
rect 13500 1943 13631 1977
rect 13034 1908 13631 1943
rect 13034 1874 13058 1908
rect 13092 1874 13126 1908
rect 13160 1874 13194 1908
rect 13228 1874 13262 1908
rect 13296 1874 13330 1908
rect 13364 1874 13398 1908
rect 13432 1874 13466 1908
rect 13500 1874 13631 1908
rect 13034 1839 13631 1874
rect 13034 1805 13058 1839
rect 13092 1805 13126 1839
rect 13160 1805 13194 1839
rect 13228 1805 13262 1839
rect 13296 1805 13330 1839
rect 13364 1805 13398 1839
rect 13432 1805 13466 1839
rect 13500 1805 13631 1839
rect 13034 1770 13631 1805
rect 13034 1736 13058 1770
rect 13092 1736 13126 1770
rect 13160 1736 13194 1770
rect 13228 1736 13262 1770
rect 13296 1736 13330 1770
rect 13364 1736 13398 1770
rect 13432 1736 13466 1770
rect 13500 1736 13631 1770
rect 13034 1701 13631 1736
rect 13034 1667 13058 1701
rect 13092 1667 13126 1701
rect 13160 1667 13194 1701
rect 13228 1667 13262 1701
rect 13296 1667 13330 1701
rect 13364 1667 13398 1701
rect 13432 1667 13466 1701
rect 13500 1667 13631 1701
rect 13034 1632 13631 1667
rect 13034 1598 13058 1632
rect 13092 1598 13126 1632
rect 13160 1598 13194 1632
rect 13228 1598 13262 1632
rect 13296 1598 13330 1632
rect 13364 1598 13398 1632
rect 13432 1598 13466 1632
rect 13500 1598 13631 1632
rect 13034 1563 13631 1598
rect 13034 1529 13058 1563
rect 13092 1529 13126 1563
rect 13160 1529 13194 1563
rect 13228 1529 13262 1563
rect 13296 1529 13330 1563
rect 13364 1529 13398 1563
rect 13432 1529 13466 1563
rect 13500 1529 13631 1563
rect 13034 1494 13631 1529
rect 13034 1426 13058 1494
rect 10619 1328 10653 1426
rect 10687 1392 10722 1426
rect 10756 1392 10791 1426
rect 10825 1392 10860 1426
rect 10894 1392 10929 1426
rect 10963 1392 10998 1426
rect 11032 1392 11067 1426
rect 11101 1392 11136 1426
rect 11170 1392 11205 1426
rect 11239 1392 11274 1426
rect 11308 1392 11343 1426
rect 11377 1392 11412 1426
rect 11446 1392 11481 1426
rect 11515 1392 11550 1426
rect 11584 1392 11619 1426
rect 11653 1392 11688 1426
rect 11722 1392 11757 1426
rect 11791 1392 11826 1426
rect 11860 1392 11895 1426
rect 11929 1392 11964 1426
rect 11998 1392 12033 1426
rect 12067 1392 12102 1426
rect 12136 1392 12171 1426
rect 12205 1392 12240 1426
rect 12274 1392 12309 1426
rect 12343 1392 12378 1426
rect 12412 1392 12447 1426
rect 12481 1392 12516 1426
rect 12550 1392 12585 1426
rect 12619 1392 12653 1426
rect 12687 1392 12721 1426
rect 12755 1392 12789 1426
rect 12823 1392 12857 1426
rect 12891 1392 12925 1426
rect 12959 1392 12993 1426
rect 13027 1392 13058 1426
rect 13231 1460 13262 1494
rect 13231 1392 13279 1460
rect 13500 1426 13631 1494
rect 13517 1392 13551 1426
rect 13585 1392 13631 1426
rect 19052 740 19154 764
rect 19086 706 19154 740
rect 19052 667 19154 706
rect 19086 633 19154 667
rect 19052 594 19154 633
rect 19086 560 19154 594
rect 19052 522 19154 560
rect 19086 488 19154 522
rect 10619 428 10653 452
rect 10619 338 10653 394
rect 19052 450 19154 488
rect 19086 416 19154 450
rect 19052 378 19154 416
rect 19086 344 19154 378
rect 10653 304 10721 328
rect 10619 294 10721 304
rect 10755 294 10790 328
rect 10824 294 10859 328
rect 10893 294 10928 328
rect 10962 294 10997 328
rect 11031 294 11066 328
rect 11100 294 11135 328
rect 11169 294 11204 328
rect 11238 294 11273 328
rect 11307 294 11342 328
rect 11376 294 11411 328
rect 11445 294 11480 328
rect 11514 294 11549 328
rect 11583 294 11618 328
rect 11652 294 11687 328
rect 11721 294 11756 328
rect 11790 294 11825 328
rect 11859 294 11894 328
rect 11928 294 11963 328
rect 11997 294 12032 328
rect 12066 294 12101 328
rect 12135 294 12170 328
rect 12204 294 12239 328
rect 12273 294 12308 328
rect 12342 294 12377 328
rect 12411 294 12446 328
rect 12480 294 12515 328
rect 12549 294 12584 328
rect 12618 294 12653 328
rect 12687 294 12722 328
rect 12756 294 12791 328
rect 12825 294 12860 328
rect 12894 294 12929 328
rect 12963 294 12998 328
rect 13032 294 13067 328
rect 10619 260 13067 294
rect 10619 248 10721 260
rect 10653 226 10721 248
rect 10755 226 10790 260
rect 10824 226 10859 260
rect 10893 226 10928 260
rect 10962 226 10997 260
rect 11031 226 11066 260
rect 11100 226 11135 260
rect 11169 226 11204 260
rect 11238 226 11273 260
rect 11307 226 11342 260
rect 11376 226 11411 260
rect 11445 226 11480 260
rect 11514 226 11549 260
rect 11583 226 11618 260
rect 11652 226 11687 260
rect 11721 226 11756 260
rect 11790 226 11825 260
rect 11859 226 11894 260
rect 11928 226 11963 260
rect 11997 226 12032 260
rect 12066 226 12101 260
rect 12135 226 12170 260
rect 12204 226 12239 260
rect 12273 226 12308 260
rect 12342 226 12377 260
rect 12411 226 12446 260
rect 12480 226 12515 260
rect 12549 226 12584 260
rect 12618 226 12653 260
rect 12687 226 12722 260
rect 12756 226 12791 260
rect 12825 226 12860 260
rect 12894 226 12929 260
rect 12963 226 12998 260
rect 13032 226 13067 260
rect 10653 214 13067 226
rect 10619 192 13067 214
rect 10619 158 10721 192
rect 10755 158 10790 192
rect 10824 158 10859 192
rect 10893 158 10928 192
rect 10962 158 10997 192
rect 11031 158 11066 192
rect 11100 158 11135 192
rect 11169 158 11204 192
rect 11238 158 11273 192
rect 11307 158 11342 192
rect 11376 158 11411 192
rect 11445 158 11480 192
rect 11514 158 11549 192
rect 11583 158 11618 192
rect 11652 158 11687 192
rect 11721 158 11756 192
rect 11790 158 11825 192
rect 11859 158 11894 192
rect 11928 158 11963 192
rect 11997 158 12032 192
rect 12066 158 12101 192
rect 12135 158 12170 192
rect 12204 158 12239 192
rect 12273 158 12308 192
rect 12342 158 12377 192
rect 12411 158 12446 192
rect 12480 158 12515 192
rect 12549 158 12584 192
rect 12618 158 12653 192
rect 12687 158 12722 192
rect 12756 158 12791 192
rect 12825 158 12860 192
rect 12894 158 12929 192
rect 12963 158 12998 192
rect 13032 158 13067 192
rect 10653 124 13067 158
rect 15073 294 15097 328
rect 19052 306 19154 344
rect 15073 260 15171 294
rect 15205 260 15240 294
rect 15274 260 15309 294
rect 15343 260 15378 294
rect 15412 260 15447 294
rect 15481 260 15516 294
rect 15550 260 15585 294
rect 15619 260 15654 294
rect 15688 260 15723 294
rect 15757 260 15792 294
rect 15826 260 15861 294
rect 15895 260 15930 294
rect 15964 260 15999 294
rect 16033 260 16068 294
rect 16102 260 16137 294
rect 16171 260 16206 294
rect 16240 260 16275 294
rect 16309 260 16344 294
rect 16378 260 16413 294
rect 16447 260 16482 294
rect 16516 260 16551 294
rect 16585 260 16620 294
rect 16654 260 16689 294
rect 16723 260 16758 294
rect 16792 260 16827 294
rect 16861 260 16896 294
rect 16930 260 16965 294
rect 16999 260 17034 294
rect 17068 260 17103 294
rect 17137 260 17172 294
rect 17206 260 17241 294
rect 17275 260 17310 294
rect 17344 260 17379 294
rect 17413 260 17448 294
rect 17482 260 17517 294
rect 17551 260 17586 294
rect 17620 260 17655 294
rect 17689 260 17724 294
rect 17758 260 17793 294
rect 17827 260 17862 294
rect 17896 260 17931 294
rect 17965 260 18000 294
rect 18034 260 18069 294
rect 18103 260 18138 294
rect 18172 260 18208 294
rect 18242 260 18278 294
rect 18312 260 18348 294
rect 18382 260 18418 294
rect 18452 260 18488 294
rect 18522 260 18558 294
rect 18592 260 18628 294
rect 18662 260 18698 294
rect 18732 260 18768 294
rect 18802 260 18838 294
rect 18872 260 18908 294
rect 18942 260 18978 294
rect 19012 272 19052 294
rect 19086 272 19154 306
rect 19012 260 19154 272
rect 15073 234 19154 260
rect 15073 226 19052 234
rect 15073 192 15171 226
rect 15205 192 15240 226
rect 15274 192 15309 226
rect 15343 192 15378 226
rect 15412 192 15447 226
rect 15481 192 15516 226
rect 15550 192 15585 226
rect 15619 192 15654 226
rect 15688 192 15723 226
rect 15757 192 15792 226
rect 15826 192 15861 226
rect 15895 192 15930 226
rect 15964 192 15999 226
rect 16033 192 16068 226
rect 16102 192 16137 226
rect 16171 192 16206 226
rect 16240 192 16275 226
rect 16309 192 16344 226
rect 16378 192 16413 226
rect 16447 192 16482 226
rect 16516 192 16551 226
rect 16585 192 16620 226
rect 16654 192 16689 226
rect 16723 192 16758 226
rect 16792 192 16827 226
rect 16861 192 16896 226
rect 16930 192 16965 226
rect 16999 192 17034 226
rect 17068 192 17103 226
rect 17137 192 17172 226
rect 17206 192 17241 226
rect 17275 192 17310 226
rect 17344 192 17379 226
rect 17413 192 17448 226
rect 17482 192 17517 226
rect 17551 192 17586 226
rect 17620 192 17655 226
rect 17689 192 17724 226
rect 17758 192 17793 226
rect 17827 192 17862 226
rect 17896 192 17931 226
rect 17965 192 18000 226
rect 18034 192 18069 226
rect 18103 192 18138 226
rect 18172 192 18208 226
rect 18242 192 18278 226
rect 18312 192 18348 226
rect 18382 192 18418 226
rect 18452 192 18488 226
rect 18522 192 18558 226
rect 18592 192 18628 226
rect 18662 192 18698 226
rect 18732 192 18768 226
rect 18802 192 18838 226
rect 18872 192 18908 226
rect 18942 192 18978 226
rect 19012 200 19052 226
rect 19086 200 19154 234
rect 19012 192 19154 200
rect 15073 124 19154 192
rect 10619 90 10721 124
rect 10755 90 10789 124
rect 10823 90 10857 124
rect 10891 90 10925 124
rect 10959 90 10993 124
rect 11027 90 11061 124
rect 11095 90 11129 124
rect 11163 90 11197 124
rect 11231 90 11265 124
rect 11299 90 11333 124
rect 11367 90 11401 124
rect 11435 90 11469 124
rect 11503 90 11537 124
rect 11571 90 11605 124
rect 11639 90 11673 124
rect 11707 90 11741 124
rect 11775 90 11809 124
rect 11843 90 11877 124
rect 11911 90 11945 124
rect 11979 90 12013 124
rect 12047 90 12081 124
rect 12115 90 12149 124
rect 12183 90 12217 124
rect 12251 90 12285 124
rect 12319 90 12353 124
rect 12387 90 12421 124
rect 12455 90 12489 124
rect 12523 90 12557 124
rect 12591 90 12625 124
rect 12659 90 12693 124
rect 12727 90 12761 124
rect 12795 90 12829 124
rect 12863 90 12897 124
rect 12931 90 12965 124
rect 12999 90 13033 124
rect 15107 90 15141 124
rect 15175 90 15209 124
rect 15243 90 15277 124
rect 15311 90 15345 124
rect 15379 90 15413 124
rect 15447 90 15481 124
rect 15515 90 15549 124
rect 15583 90 15617 124
rect 15651 90 15685 124
rect 15719 90 15753 124
rect 15787 90 15821 124
rect 15855 90 15889 124
rect 15923 90 15957 124
rect 15991 90 16025 124
rect 16059 90 16093 124
rect 16127 90 16161 124
rect 16195 90 16229 124
rect 16263 90 16297 124
rect 16331 90 16365 124
rect 16399 90 16433 124
rect 16467 90 16501 124
rect 16535 90 16569 124
rect 16603 90 16637 124
rect 16671 90 16705 124
rect 16739 90 16773 124
rect 16807 90 16841 124
rect 16875 90 16909 124
rect 16943 90 16977 124
rect 17011 90 17045 124
rect 17079 90 17113 124
rect 17147 90 17181 124
rect 17215 90 17249 124
rect 17283 90 17317 124
rect 17351 90 17385 124
rect 17419 90 17453 124
rect 17487 90 17521 124
rect 17555 90 17589 124
rect 17623 90 17657 124
rect 17691 90 17725 124
rect 17759 90 17793 124
rect 17827 90 17861 124
rect 17895 90 17929 124
rect 17963 90 17997 124
rect 18031 90 18065 124
rect 18099 90 18133 124
rect 18167 90 18201 124
rect 18235 90 18269 124
rect 18303 90 18337 124
rect 18371 90 18405 124
rect 18439 90 18473 124
rect 18507 90 18541 124
rect 18575 90 18609 124
rect 18643 90 18677 124
rect 18711 90 18745 124
rect 18779 90 18813 124
rect 18847 90 18881 124
rect 18915 90 18949 124
rect 18983 90 19018 124
rect 19052 90 19154 124
rect 18872 64 19154 90
<< mvnsubdiff >>
rect -25 6906 -1 6940
rect 33 6906 68 6940
rect 102 6906 137 6940
rect 171 6906 206 6940
rect 240 6906 275 6940
rect 309 6906 344 6940
rect 378 6906 413 6940
rect 447 6906 482 6940
rect 516 6906 551 6940
rect 585 6906 620 6940
rect 654 6906 689 6940
rect 723 6906 758 6940
rect 792 6906 827 6940
rect 861 6906 896 6940
rect 930 6906 965 6940
rect 999 6906 1034 6940
rect 1068 6906 1103 6940
rect 1137 6906 1172 6940
rect 1206 6906 1241 6940
rect 1275 6906 1310 6940
rect 1344 6906 1379 6940
rect 1413 6906 1448 6940
rect 1482 6906 1517 6940
rect 1551 6906 1586 6940
rect 1620 6906 1655 6940
rect 1689 6906 1724 6940
rect 1758 6906 1793 6940
rect 1827 6906 1862 6940
rect -25 6872 1862 6906
rect -25 6838 -1 6872
rect 33 6838 68 6872
rect 102 6838 137 6872
rect 171 6838 206 6872
rect 240 6838 275 6872
rect 309 6838 344 6872
rect 378 6838 413 6872
rect 447 6838 482 6872
rect 516 6838 551 6872
rect 585 6838 620 6872
rect 654 6838 689 6872
rect 723 6838 758 6872
rect 792 6838 827 6872
rect 861 6838 896 6872
rect 930 6838 965 6872
rect 999 6838 1034 6872
rect 1068 6838 1103 6872
rect 1137 6838 1172 6872
rect 1206 6838 1241 6872
rect 1275 6838 1310 6872
rect 1344 6838 1379 6872
rect 1413 6838 1448 6872
rect 1482 6838 1517 6872
rect 1551 6838 1586 6872
rect 1620 6838 1655 6872
rect 1689 6838 1724 6872
rect 1758 6838 1793 6872
rect 1827 6838 1862 6872
rect -25 6804 1862 6838
rect -25 6770 -1 6804
rect 33 6770 68 6804
rect 102 6770 137 6804
rect 171 6770 206 6804
rect 240 6770 275 6804
rect 309 6770 344 6804
rect 378 6770 413 6804
rect 447 6770 482 6804
rect 516 6770 551 6804
rect 585 6770 620 6804
rect 654 6770 689 6804
rect 723 6770 758 6804
rect 792 6770 827 6804
rect 861 6770 896 6804
rect 930 6770 965 6804
rect 999 6770 1034 6804
rect 1068 6770 1103 6804
rect 1137 6770 1172 6804
rect 1206 6770 1241 6804
rect 1275 6770 1310 6804
rect 1344 6770 1379 6804
rect 1413 6770 1448 6804
rect 1482 6770 1517 6804
rect 1551 6770 1586 6804
rect 1620 6770 1655 6804
rect 1689 6770 1724 6804
rect 1758 6770 1793 6804
rect 1827 6770 1862 6804
rect 10056 6906 10090 6940
rect 10124 6906 10158 6940
rect 10192 6906 10226 6940
rect 10260 6906 10294 6940
rect 10328 6906 10362 6940
rect 10396 6906 10430 6940
rect 10464 6906 10498 6940
rect 10532 6906 10566 6940
rect 10600 6906 10634 6940
rect 10668 6906 10702 6940
rect 10736 6906 10770 6940
rect 10804 6906 10838 6940
rect 10872 6906 10906 6940
rect 10940 6906 10974 6940
rect 11008 6906 11042 6940
rect 11076 6906 11110 6940
rect 11144 6906 11178 6940
rect 11212 6906 11246 6940
rect 11280 6906 11314 6940
rect 11348 6906 11382 6940
rect 11416 6906 11450 6940
rect 11484 6906 11518 6940
rect 11552 6906 11586 6940
rect 11620 6906 11654 6940
rect 11688 6906 11722 6940
rect 11756 6906 11790 6940
rect 11824 6906 11858 6940
rect 11892 6906 11926 6940
rect 11960 6906 11994 6940
rect 12028 6906 12062 6940
rect 12096 6906 12130 6940
rect 12164 6906 12198 6940
rect 12232 6906 12266 6940
rect 12300 6906 12334 6940
rect 12368 6906 12402 6940
rect 12436 6906 12471 6940
rect 12505 6906 12540 6940
rect 12574 6906 12609 6940
rect 12643 6906 12678 6940
rect 12712 6906 12747 6940
rect 12781 6906 12816 6940
rect 12850 6906 12885 6940
rect 12919 6906 12954 6940
rect 12988 6906 13023 6940
rect 13057 6906 13092 6940
rect 13126 6906 13161 6940
rect 13195 6906 13230 6940
rect 13264 6906 13299 6940
rect 13333 6906 13367 6940
rect 10056 6872 13367 6906
rect 10056 6838 10091 6872
rect 10125 6838 10160 6872
rect 10194 6838 10229 6872
rect 10263 6838 10298 6872
rect 10332 6838 10367 6872
rect 10401 6838 10436 6872
rect 10470 6838 10505 6872
rect 10539 6838 10574 6872
rect 10608 6838 10643 6872
rect 10677 6838 10712 6872
rect 10746 6838 10781 6872
rect 10815 6838 10850 6872
rect 10884 6838 10919 6872
rect 10953 6838 10988 6872
rect 11022 6838 11057 6872
rect 11091 6838 11126 6872
rect 11160 6838 11195 6872
rect 11229 6838 11264 6872
rect 11298 6838 11333 6872
rect 11367 6838 11402 6872
rect 11436 6838 11471 6872
rect 11505 6838 11540 6872
rect 11574 6838 11609 6872
rect 11643 6838 11678 6872
rect 11712 6838 11747 6872
rect 11781 6838 11816 6872
rect 11850 6838 11885 6872
rect 11919 6838 11954 6872
rect 11988 6838 12023 6872
rect 12057 6838 12092 6872
rect 12126 6838 12161 6872
rect 12195 6838 12230 6872
rect 12264 6838 12299 6872
rect 12333 6838 12368 6872
rect 12402 6838 12437 6872
rect 12471 6838 12506 6872
rect 12540 6838 12575 6872
rect 12609 6838 12644 6872
rect 12678 6838 12713 6872
rect 12747 6838 12782 6872
rect 12816 6838 12851 6872
rect 12885 6838 12920 6872
rect 12954 6838 12989 6872
rect 13023 6838 13058 6872
rect 13092 6838 13127 6872
rect 13161 6838 13196 6872
rect 13230 6838 13265 6872
rect 13299 6838 13367 6872
rect 10056 6804 13265 6838
rect 10056 6770 10091 6804
rect 10125 6770 10160 6804
rect 10194 6770 10229 6804
rect 10263 6770 10298 6804
rect 10332 6770 10367 6804
rect 10401 6770 10436 6804
rect 10470 6770 10505 6804
rect 10539 6770 10574 6804
rect 10608 6770 10643 6804
rect 10677 6770 10712 6804
rect 10746 6770 10781 6804
rect 10815 6770 10850 6804
rect 10884 6770 10919 6804
rect 10953 6770 10988 6804
rect 11022 6770 11057 6804
rect 11091 6770 11126 6804
rect 11160 6770 11195 6804
rect 11229 6770 11264 6804
rect 11298 6770 11333 6804
rect 11367 6770 11402 6804
rect 11436 6770 11471 6804
rect 11505 6770 11540 6804
rect 11574 6770 11609 6804
rect 11643 6770 11678 6804
rect 11712 6770 11747 6804
rect 11781 6770 11816 6804
rect 11850 6770 11885 6804
rect 11919 6770 11954 6804
rect 11988 6770 12023 6804
rect 12057 6770 12092 6804
rect 12126 6770 12161 6804
rect 12195 6770 12230 6804
rect 12264 6770 12299 6804
rect 12333 6770 12368 6804
rect 12402 6770 12437 6804
rect 12471 6770 12506 6804
rect 12540 6770 12575 6804
rect 12609 6770 12644 6804
rect 12678 6770 12713 6804
rect 12747 6770 12782 6804
rect 12816 6770 12851 6804
rect 12885 6770 12920 6804
rect 12954 6770 12989 6804
rect 13023 6770 13058 6804
rect 13092 6770 13127 6804
rect 13161 6770 13197 6804
rect 2533 6751 13197 6770
rect 3340 6728 5568 6751
rect 3340 6694 3373 6728
rect 3407 6694 3441 6728
rect 3475 6694 3509 6728
rect 3543 6694 3577 6728
rect 3611 6694 3645 6728
rect 3679 6694 3713 6728
rect 3747 6694 3781 6728
rect 3815 6694 3849 6728
rect 3883 6694 3917 6728
rect 3951 6694 3985 6728
rect 4019 6694 4053 6728
rect 4087 6694 4121 6728
rect 4155 6694 4189 6728
rect 4223 6694 4257 6728
rect 4291 6694 4325 6728
rect 4359 6694 4393 6728
rect 4427 6694 4461 6728
rect 4495 6694 4529 6728
rect 4563 6694 4597 6728
rect 4631 6694 4665 6728
rect 4699 6694 4733 6728
rect 4767 6694 4801 6728
rect 4835 6694 4869 6728
rect 4903 6694 4937 6728
rect 4971 6694 5005 6728
rect 5039 6694 5073 6728
rect 5107 6695 5568 6728
rect 5107 6694 5180 6695
rect 3340 6661 5180 6694
rect 5214 6661 5248 6695
rect 5282 6661 5316 6695
rect 5350 6661 5384 6695
rect 5418 6661 5452 6695
rect 5486 6661 5520 6695
rect 5554 6661 5568 6695
rect 3340 6658 5568 6661
rect 3340 6624 3373 6658
rect 3407 6624 3441 6658
rect 3475 6624 3509 6658
rect 3543 6624 3577 6658
rect 3611 6624 3645 6658
rect 3679 6624 3713 6658
rect 3747 6624 3781 6658
rect 3815 6624 3849 6658
rect 3883 6624 3917 6658
rect 3951 6624 3985 6658
rect 4019 6624 4053 6658
rect 4087 6624 4121 6658
rect 4155 6624 4189 6658
rect 4223 6624 4257 6658
rect 4291 6624 4325 6658
rect 4359 6624 4393 6658
rect 4427 6624 4461 6658
rect 4495 6624 4529 6658
rect 4563 6624 4597 6658
rect 4631 6624 4665 6658
rect 4699 6624 4733 6658
rect 4767 6624 4801 6658
rect 4835 6624 4869 6658
rect 4903 6624 4937 6658
rect 4971 6624 5005 6658
rect 5039 6624 5073 6658
rect 5107 6625 5568 6658
rect 5107 6624 5180 6625
rect 3340 6591 5180 6624
rect 5214 6591 5248 6625
rect 5282 6591 5316 6625
rect 5350 6591 5384 6625
rect 5418 6591 5452 6625
rect 5486 6591 5520 6625
rect 5554 6591 5568 6625
rect 6781 6736 6815 6751
rect 6781 6663 6815 6702
rect 3340 6588 5568 6591
rect 3340 6554 3373 6588
rect 3407 6554 3441 6588
rect 3475 6554 3509 6588
rect 3543 6554 3577 6588
rect 3611 6554 3645 6588
rect 3679 6554 3713 6588
rect 3747 6554 3781 6588
rect 3815 6554 3849 6588
rect 3883 6554 3917 6588
rect 3951 6554 3985 6588
rect 4019 6554 4053 6588
rect 4087 6554 4121 6588
rect 4155 6554 4189 6588
rect 4223 6554 4257 6588
rect 4291 6554 4325 6588
rect 4359 6554 4393 6588
rect 4427 6554 4461 6588
rect 4495 6554 4529 6588
rect 4563 6554 4597 6588
rect 4631 6554 4665 6588
rect 4699 6554 4733 6588
rect 4767 6554 4801 6588
rect 4835 6554 4869 6588
rect 4903 6554 4937 6588
rect 4971 6554 5005 6588
rect 5039 6554 5073 6588
rect 5107 6556 5568 6588
rect 5107 6554 5180 6556
rect 3340 6522 5180 6554
rect 5214 6522 5248 6556
rect 5282 6522 5316 6556
rect 5350 6522 5384 6556
rect 5418 6522 5452 6556
rect 5486 6522 5520 6556
rect 5554 6522 5568 6556
rect 3340 6518 5568 6522
rect 3340 6484 3373 6518
rect 3407 6484 3441 6518
rect 3475 6484 3509 6518
rect 3543 6484 3577 6518
rect 3611 6484 3645 6518
rect 3679 6484 3713 6518
rect 3747 6484 3781 6518
rect 3815 6484 3849 6518
rect 3883 6484 3917 6518
rect 3951 6484 3985 6518
rect 4019 6484 4053 6518
rect 4087 6484 4121 6518
rect 4155 6484 4189 6518
rect 4223 6484 4257 6518
rect 4291 6484 4325 6518
rect 4359 6484 4393 6518
rect 4427 6484 4461 6518
rect 4495 6484 4529 6518
rect 4563 6484 4597 6518
rect 4631 6484 4665 6518
rect 4699 6484 4733 6518
rect 4767 6484 4801 6518
rect 4835 6484 4869 6518
rect 4903 6484 4937 6518
rect 4971 6484 5005 6518
rect 5039 6484 5073 6518
rect 5107 6487 5568 6518
rect 5107 6484 5180 6487
rect 3340 6453 5180 6484
rect 5214 6453 5248 6487
rect 5282 6453 5316 6487
rect 5350 6453 5384 6487
rect 5418 6453 5452 6487
rect 5486 6453 5520 6487
rect 5554 6453 5568 6487
rect 3340 6448 5568 6453
rect 3340 6414 3373 6448
rect 3407 6414 3441 6448
rect 3475 6414 3509 6448
rect 3543 6414 3577 6448
rect 3611 6414 3645 6448
rect 3679 6414 3713 6448
rect 3747 6414 3781 6448
rect 3815 6414 3849 6448
rect 3883 6414 3917 6448
rect 3951 6414 3985 6448
rect 4019 6414 4053 6448
rect 4087 6414 4121 6448
rect 4155 6414 4189 6448
rect 4223 6414 4257 6448
rect 4291 6414 4325 6448
rect 4359 6414 4393 6448
rect 4427 6414 4461 6448
rect 4495 6414 4529 6448
rect 4563 6414 4597 6448
rect 4631 6414 4665 6448
rect 4699 6414 4733 6448
rect 4767 6414 4801 6448
rect 4835 6414 4869 6448
rect 4903 6414 4937 6448
rect 4971 6414 5005 6448
rect 5039 6414 5073 6448
rect 5107 6418 5568 6448
rect 6781 6591 6815 6629
rect 6781 6519 6815 6557
rect 6781 6448 6815 6485
rect 9283 6720 13197 6751
rect 9283 6448 9317 6720
rect 13159 6482 13197 6720
rect 5107 6414 5180 6418
rect 3340 6384 5180 6414
rect 5214 6384 5248 6418
rect 5282 6384 5316 6418
rect 5350 6384 5384 6418
rect 5418 6384 5452 6418
rect 5486 6384 5520 6418
rect 5554 6384 5568 6418
rect 6781 6414 6825 6448
rect 6859 6414 6893 6448
rect 6927 6414 6961 6448
rect 6995 6414 7029 6448
rect 7063 6414 7097 6448
rect 7131 6414 7165 6448
rect 7199 6414 7233 6448
rect 7267 6414 7301 6448
rect 7335 6414 7369 6448
rect 7403 6414 7437 6448
rect 7471 6414 7505 6448
rect 7539 6414 7573 6448
rect 7607 6414 7641 6448
rect 7675 6414 7709 6448
rect 7743 6414 7777 6448
rect 7811 6414 7845 6448
rect 7879 6414 7913 6448
rect 7947 6414 7981 6448
rect 8015 6414 8049 6448
rect 8083 6414 8117 6448
rect 8151 6414 8185 6448
rect 8219 6414 8253 6448
rect 8287 6414 8321 6448
rect 8355 6414 8389 6448
rect 8423 6414 8457 6448
rect 8491 6414 8525 6448
rect 8559 6414 8593 6448
rect 8627 6414 8661 6448
rect 8695 6414 8729 6448
rect 8763 6414 8797 6448
rect 8831 6414 8865 6448
rect 8899 6414 8933 6448
rect 8967 6414 9001 6448
rect 9035 6414 9069 6448
rect 9103 6414 9137 6448
rect 9171 6414 9205 6448
rect 9239 6414 9273 6448
rect 9307 6414 9317 6448
rect 9851 6448 13197 6482
rect 9851 6414 9886 6448
rect 9920 6414 9955 6448
rect 9989 6414 10024 6448
rect 10058 6414 10093 6448
rect 10127 6414 10162 6448
rect 10196 6414 10231 6448
rect 10265 6414 10300 6448
rect 10334 6414 10369 6448
rect 10403 6414 10438 6448
rect 10472 6414 10507 6448
rect 10541 6414 10576 6448
rect 10610 6414 10645 6448
rect 10679 6414 10714 6448
rect 10748 6414 10783 6448
rect 10817 6414 10852 6448
rect 10886 6414 10921 6448
rect 10955 6414 10990 6448
rect 11024 6414 11059 6448
rect 11093 6414 11128 6448
rect 11162 6414 11197 6448
rect 11231 6414 11266 6448
rect 11300 6414 11335 6448
rect 11369 6414 11404 6448
rect 11438 6414 11473 6448
rect 11507 6414 11542 6448
rect 11576 6414 11611 6448
rect 11645 6414 11680 6448
rect 11714 6414 11749 6448
rect 11783 6414 11818 6448
rect 11852 6414 11887 6448
rect 11921 6414 11956 6448
rect 11990 6414 12025 6448
rect 12059 6414 12094 6448
rect 12128 6414 12163 6448
rect 12197 6414 12232 6448
rect 12266 6414 12301 6448
rect 12335 6414 12370 6448
rect 12404 6414 12439 6448
rect 12473 6414 12508 6448
rect 12542 6414 12577 6448
rect 12611 6414 12646 6448
rect 12680 6414 12715 6448
rect 12749 6414 12784 6448
rect 12818 6414 12853 6448
rect 12887 6414 12922 6448
rect 12956 6414 12991 6448
rect 13025 6414 13060 6448
rect 13094 6414 13129 6448
rect 13163 6414 13197 6448
rect 3340 6378 5568 6384
rect 3340 6344 3373 6378
rect 3407 6344 3441 6378
rect 3475 6344 3509 6378
rect 3543 6344 3577 6378
rect 3611 6344 3645 6378
rect 3679 6344 3713 6378
rect 3747 6344 3781 6378
rect 3815 6344 3849 6378
rect 3883 6344 3917 6378
rect 3951 6344 3985 6378
rect 4019 6344 4053 6378
rect 4087 6344 4121 6378
rect 4155 6344 4189 6378
rect 4223 6344 4257 6378
rect 4291 6344 4325 6378
rect 4359 6344 4393 6378
rect 4427 6344 4461 6378
rect 4495 6344 4529 6378
rect 4563 6344 4597 6378
rect 4631 6344 4665 6378
rect 4699 6344 4733 6378
rect 4767 6344 4801 6378
rect 4835 6344 4869 6378
rect 4903 6344 4937 6378
rect 4971 6344 5005 6378
rect 5039 6344 5073 6378
rect 5107 6349 5568 6378
rect 5107 6344 5180 6349
rect 3340 6315 5180 6344
rect 5214 6315 5248 6349
rect 5282 6315 5316 6349
rect 5350 6315 5384 6349
rect 5418 6315 5452 6349
rect 5486 6315 5520 6349
rect 5554 6315 5568 6349
rect 3340 6308 5568 6315
rect 3340 6274 3373 6308
rect 3407 6274 3441 6308
rect 3475 6274 3509 6308
rect 3543 6274 3577 6308
rect 3611 6274 3645 6308
rect 3679 6274 3713 6308
rect 3747 6274 3781 6308
rect 3815 6274 3849 6308
rect 3883 6274 3917 6308
rect 3951 6274 3985 6308
rect 4019 6274 4053 6308
rect 4087 6274 4121 6308
rect 4155 6274 4189 6308
rect 4223 6274 4257 6308
rect 4291 6274 4325 6308
rect 4359 6274 4393 6308
rect 4427 6274 4461 6308
rect 4495 6274 4529 6308
rect 4563 6274 4597 6308
rect 4631 6274 4665 6308
rect 4699 6274 4733 6308
rect 4767 6274 4801 6308
rect 4835 6274 4869 6308
rect 4903 6274 4937 6308
rect 4971 6274 5005 6308
rect 5039 6274 5073 6308
rect 5107 6274 5568 6308
rect 3340 6242 5568 6274
rect 3340 6238 6781 6242
rect 3340 6204 3373 6238
rect 3407 6204 3441 6238
rect 3475 6204 3509 6238
rect 3543 6204 3577 6238
rect 3611 6204 3645 6238
rect 3679 6204 3713 6238
rect 3747 6204 3781 6238
rect 3815 6204 3849 6238
rect 3883 6204 3917 6238
rect 3951 6204 3985 6238
rect 4019 6204 4053 6238
rect 4087 6204 4121 6238
rect 4155 6204 4189 6238
rect 4223 6204 4257 6238
rect 4291 6204 4325 6238
rect 4359 6204 4393 6238
rect 4427 6204 4461 6238
rect 4495 6204 4529 6238
rect 4563 6204 4597 6238
rect 4631 6204 4665 6238
rect 4699 6204 4733 6238
rect 4767 6204 4801 6238
rect 4835 6204 4869 6238
rect 4903 6204 4937 6238
rect 4971 6204 5005 6238
rect 5039 6204 5073 6238
rect 5107 6218 6781 6238
rect 5107 6204 5155 6218
rect 3340 6184 5155 6204
rect 5189 6184 5223 6218
rect 5257 6184 5291 6218
rect 5325 6184 5359 6218
rect 5393 6184 5427 6218
rect 5461 6184 5495 6218
rect 5529 6184 5563 6218
rect 5597 6184 5631 6218
rect 5665 6184 5699 6218
rect 5733 6184 5767 6218
rect 5801 6184 5835 6218
rect 5869 6184 5903 6218
rect 5937 6184 5971 6218
rect 6005 6184 6040 6218
rect 6074 6184 6108 6218
rect 6142 6184 6176 6218
rect 6210 6184 6244 6218
rect 6278 6184 6312 6218
rect 6346 6184 6380 6218
rect 6414 6184 6448 6218
rect 6482 6184 6516 6218
rect 6550 6184 6584 6218
rect 6618 6184 6652 6218
rect 6686 6184 6720 6218
rect 6754 6184 6781 6218
rect 3340 6168 6781 6184
rect 3340 6134 3373 6168
rect 3407 6134 3441 6168
rect 3475 6134 3509 6168
rect 3543 6134 3577 6168
rect 3611 6134 3645 6168
rect 3679 6134 3713 6168
rect 3747 6134 3781 6168
rect 3815 6134 3849 6168
rect 3883 6134 3917 6168
rect 3951 6134 3985 6168
rect 4019 6134 4053 6168
rect 4087 6134 4121 6168
rect 4155 6134 4189 6168
rect 4223 6134 4257 6168
rect 4291 6134 4325 6168
rect 4359 6134 4393 6168
rect 4427 6134 4461 6168
rect 4495 6134 4529 6168
rect 4563 6134 4597 6168
rect 4631 6134 4665 6168
rect 4699 6134 4733 6168
rect 4767 6134 4801 6168
rect 4835 6134 4869 6168
rect 4903 6134 4937 6168
rect 4971 6134 5005 6168
rect 5039 6134 5073 6168
rect 5107 6149 6781 6168
rect 5107 6148 6040 6149
rect 5107 6134 5155 6148
rect 3340 6114 5155 6134
rect 5189 6114 5223 6148
rect 5257 6114 5291 6148
rect 5325 6114 5359 6148
rect 5393 6114 5427 6148
rect 5461 6114 5495 6148
rect 5529 6114 5563 6148
rect 5597 6114 5631 6148
rect 5665 6114 5699 6148
rect 5733 6114 5767 6148
rect 5801 6114 5835 6148
rect 5869 6114 5903 6148
rect 5937 6114 5971 6148
rect 6005 6115 6040 6148
rect 6074 6115 6108 6149
rect 6142 6115 6176 6149
rect 6210 6115 6244 6149
rect 6278 6115 6312 6149
rect 6346 6115 6380 6149
rect 6414 6115 6448 6149
rect 6482 6115 6516 6149
rect 6550 6115 6584 6149
rect 6618 6115 6652 6149
rect 6686 6115 6720 6149
rect 6754 6115 6781 6149
rect 6005 6114 6781 6115
rect 3340 6098 6781 6114
rect 3340 6064 3373 6098
rect 3407 6064 3441 6098
rect 3475 6064 3509 6098
rect 3543 6064 3577 6098
rect 3611 6064 3645 6098
rect 3679 6064 3713 6098
rect 3747 6064 3781 6098
rect 3815 6064 3849 6098
rect 3883 6064 3917 6098
rect 3951 6064 3985 6098
rect 4019 6064 4053 6098
rect 4087 6064 4121 6098
rect 4155 6064 4189 6098
rect 4223 6064 4257 6098
rect 4291 6064 4325 6098
rect 4359 6064 4393 6098
rect 4427 6064 4461 6098
rect 4495 6064 4529 6098
rect 4563 6064 4597 6098
rect 4631 6064 4665 6098
rect 4699 6064 4733 6098
rect 4767 6064 4801 6098
rect 4835 6064 4869 6098
rect 4903 6064 4937 6098
rect 4971 6064 5005 6098
rect 5039 6064 5073 6098
rect 5107 6080 6781 6098
rect 5107 6078 6040 6080
rect 5107 6064 5155 6078
rect 3340 6044 5155 6064
rect 5189 6044 5223 6078
rect 5257 6044 5291 6078
rect 5325 6044 5359 6078
rect 5393 6044 5427 6078
rect 5461 6044 5495 6078
rect 5529 6044 5563 6078
rect 5597 6044 5631 6078
rect 5665 6044 5699 6078
rect 5733 6044 5767 6078
rect 5801 6044 5835 6078
rect 5869 6044 5903 6078
rect 5937 6044 5971 6078
rect 6005 6046 6040 6078
rect 6074 6046 6108 6080
rect 6142 6046 6176 6080
rect 6210 6046 6244 6080
rect 6278 6046 6312 6080
rect 6346 6046 6380 6080
rect 6414 6046 6448 6080
rect 6482 6046 6516 6080
rect 6550 6046 6584 6080
rect 6618 6046 6652 6080
rect 6686 6046 6720 6080
rect 6754 6071 6781 6080
rect 6754 6046 6825 6071
rect 6005 6044 6825 6046
rect 3340 6037 6825 6044
rect 6859 6037 6893 6071
rect 6927 6037 6961 6071
rect 6995 6037 7029 6071
rect 7063 6037 7097 6071
rect 7131 6037 7165 6071
rect 7199 6037 7233 6071
rect 7267 6037 7301 6071
rect 7335 6037 7369 6071
rect 7403 6037 7437 6071
rect 7471 6037 7505 6071
rect 7539 6037 7573 6071
rect 7607 6037 7641 6071
rect 7675 6037 7709 6071
rect 7743 6037 7777 6071
rect 7811 6037 7845 6071
rect 7879 6037 7913 6071
rect 7947 6037 7981 6071
rect 8015 6037 8049 6071
rect 8083 6037 8117 6071
rect 8151 6037 8185 6071
rect 8219 6037 8253 6071
rect 8287 6037 8321 6071
rect 8355 6037 8389 6071
rect 8423 6037 8457 6071
rect 8491 6037 8525 6071
rect 8559 6037 8593 6071
rect 8627 6037 8661 6071
rect 8695 6037 8729 6071
rect 8763 6037 8797 6071
rect 8831 6037 8865 6071
rect 8899 6037 8933 6071
rect 8967 6037 9001 6071
rect 9035 6037 9069 6071
rect 9103 6037 9137 6071
rect 9171 6037 9205 6071
rect 9239 6037 9273 6071
rect 9307 6037 9341 6071
rect 9375 6037 9409 6071
rect 9443 6037 9477 6071
rect 9511 6037 9545 6071
rect 9579 6037 9613 6071
rect 9647 6037 9681 6071
rect 9715 6037 9749 6071
rect 9783 6037 9817 6071
rect 9851 6037 9886 6071
rect 9920 6037 9955 6071
rect 9989 6037 10024 6071
rect 10058 6037 10093 6071
rect 10127 6037 10162 6071
rect 10196 6037 10231 6071
rect 10265 6037 10300 6071
rect 10334 6037 10369 6071
rect 10403 6037 10438 6071
rect 10472 6037 10507 6071
rect 10541 6037 10576 6071
rect 10610 6037 10645 6071
rect 10679 6037 10714 6071
rect 10748 6037 10783 6071
rect 10817 6037 10852 6071
rect 10886 6037 10921 6071
rect 10955 6037 10990 6071
rect 11024 6037 11059 6071
rect 11093 6037 11128 6071
rect 11162 6037 11197 6071
rect 11231 6037 11266 6071
rect 11300 6037 11335 6071
rect 11369 6037 11404 6071
rect 11438 6037 11473 6071
rect 11507 6037 11542 6071
rect 11576 6037 11611 6071
rect 11645 6037 11680 6071
rect 11714 6037 11749 6071
rect 11783 6037 11818 6071
rect 11852 6037 11887 6071
rect 11921 6037 11956 6071
rect 11990 6037 12025 6071
rect 12059 6037 12094 6071
rect 12128 6037 12163 6071
rect 12197 6037 12232 6071
rect 12266 6037 12301 6071
rect 12335 6037 12370 6071
rect 12404 6037 12439 6071
rect 12473 6037 12508 6071
rect 12542 6037 12577 6071
rect 12611 6037 12646 6071
rect 12680 6037 12715 6071
rect 12749 6037 12784 6071
rect 12818 6037 12853 6071
rect 12887 6037 12922 6071
rect 12956 6037 12991 6071
rect 13025 6037 13060 6071
rect 13094 6037 13129 6071
rect 13163 6037 13197 6071
rect 3340 6028 6781 6037
rect 3340 5994 3373 6028
rect 3407 5994 3441 6028
rect 3475 5994 3509 6028
rect 3543 5994 3577 6028
rect 3611 5994 3645 6028
rect 3679 5994 3713 6028
rect 3747 5994 3781 6028
rect 3815 5994 3849 6028
rect 3883 5994 3917 6028
rect 3951 5994 3985 6028
rect 4019 5994 4053 6028
rect 4087 5994 4121 6028
rect 4155 5994 4189 6028
rect 4223 5994 4257 6028
rect 4291 5994 4325 6028
rect 4359 5994 4393 6028
rect 4427 5994 4461 6028
rect 4495 5994 4529 6028
rect 4563 5994 4597 6028
rect 4631 5994 4665 6028
rect 4699 5994 4733 6028
rect 4767 5994 4801 6028
rect 4835 5994 4869 6028
rect 4903 5994 4937 6028
rect 4971 5994 5005 6028
rect 5039 5994 5073 6028
rect 5107 6011 6781 6028
rect 5107 6008 6040 6011
rect 5107 5994 5155 6008
rect 3340 5974 5155 5994
rect 5189 5974 5223 6008
rect 5257 5974 5291 6008
rect 5325 5974 5359 6008
rect 5393 5974 5427 6008
rect 5461 5974 5495 6008
rect 5529 5974 5563 6008
rect 5597 5974 5631 6008
rect 5665 5974 5699 6008
rect 5733 5974 5767 6008
rect 5801 5974 5835 6008
rect 5869 5974 5903 6008
rect 5937 5974 5971 6008
rect 6005 5977 6040 6008
rect 6074 5977 6108 6011
rect 6142 5977 6176 6011
rect 6210 5977 6244 6011
rect 6278 5977 6312 6011
rect 6346 5977 6380 6011
rect 6414 5977 6448 6011
rect 6482 5977 6516 6011
rect 6550 5977 6584 6011
rect 6618 5977 6652 6011
rect 6686 5977 6720 6011
rect 6754 5977 6781 6011
rect 6005 5974 6781 5977
rect 3340 5958 6781 5974
rect 3340 5924 3373 5958
rect 3407 5924 3441 5958
rect 3475 5924 3509 5958
rect 3543 5924 3577 5958
rect 3611 5924 3645 5958
rect 3679 5924 3713 5958
rect 3747 5924 3781 5958
rect 3815 5924 3849 5958
rect 3883 5924 3917 5958
rect 3951 5924 3985 5958
rect 4019 5924 4053 5958
rect 4087 5924 4121 5958
rect 4155 5924 4189 5958
rect 4223 5924 4257 5958
rect 4291 5924 4325 5958
rect 4359 5924 4393 5958
rect 4427 5924 4461 5958
rect 4495 5924 4529 5958
rect 4563 5924 4597 5958
rect 4631 5924 4665 5958
rect 4699 5924 4733 5958
rect 4767 5924 4801 5958
rect 4835 5924 4869 5958
rect 4903 5924 4937 5958
rect 4971 5924 5005 5958
rect 5039 5924 5073 5958
rect 5107 5942 6781 5958
rect 5107 5938 6040 5942
rect 5107 5924 5155 5938
rect 3340 5904 5155 5924
rect 5189 5904 5223 5938
rect 5257 5904 5291 5938
rect 5325 5904 5359 5938
rect 5393 5904 5427 5938
rect 5461 5904 5495 5938
rect 5529 5904 5563 5938
rect 5597 5904 5631 5938
rect 5665 5904 5699 5938
rect 5733 5904 5767 5938
rect 5801 5904 5835 5938
rect 5869 5904 5903 5938
rect 5937 5904 5971 5938
rect 6005 5908 6040 5938
rect 6074 5908 6108 5942
rect 6142 5908 6176 5942
rect 6210 5908 6244 5942
rect 6278 5908 6312 5942
rect 6346 5908 6380 5942
rect 6414 5908 6448 5942
rect 6482 5908 6516 5942
rect 6550 5908 6584 5942
rect 6618 5908 6652 5942
rect 6686 5908 6720 5942
rect 6754 5908 6781 5942
rect 6005 5904 6781 5908
rect 3340 5888 6781 5904
rect 3340 5854 3373 5888
rect 3407 5854 3441 5888
rect 3475 5854 3509 5888
rect 3543 5854 3577 5888
rect 3611 5854 3645 5888
rect 3679 5854 3713 5888
rect 3747 5854 3781 5888
rect 3815 5854 3849 5888
rect 3883 5854 3917 5888
rect 3951 5854 3985 5888
rect 4019 5854 4053 5888
rect 4087 5854 4121 5888
rect 4155 5854 4189 5888
rect 4223 5854 4257 5888
rect 4291 5854 4325 5888
rect 4359 5854 4393 5888
rect 4427 5854 4461 5888
rect 4495 5854 4529 5888
rect 4563 5854 4597 5888
rect 4631 5854 4665 5888
rect 4699 5854 4733 5888
rect 4767 5854 4801 5888
rect 4835 5854 4869 5888
rect 4903 5854 4937 5888
rect 4971 5854 5005 5888
rect 5039 5854 5073 5888
rect 5107 5873 6781 5888
rect 5107 5868 6040 5873
rect 5107 5854 5155 5868
rect 3340 5834 5155 5854
rect 5189 5834 5223 5868
rect 5257 5834 5291 5868
rect 5325 5834 5359 5868
rect 5393 5834 5427 5868
rect 5461 5834 5495 5868
rect 5529 5834 5563 5868
rect 5597 5834 5631 5868
rect 5665 5834 5699 5868
rect 5733 5834 5767 5868
rect 5801 5834 5835 5868
rect 5869 5834 5903 5868
rect 5937 5834 5971 5868
rect 6005 5839 6040 5868
rect 6074 5839 6108 5873
rect 6142 5839 6176 5873
rect 6210 5839 6244 5873
rect 6278 5839 6312 5873
rect 6346 5839 6380 5873
rect 6414 5839 6448 5873
rect 6482 5839 6516 5873
rect 6550 5839 6584 5873
rect 6618 5839 6652 5873
rect 6686 5839 6720 5873
rect 6754 5839 6781 5873
rect 6005 5834 6781 5839
rect 3340 5818 6781 5834
rect 3340 5784 3373 5818
rect 3407 5784 3441 5818
rect 3475 5784 3509 5818
rect 3543 5784 3577 5818
rect 3611 5784 3645 5818
rect 3679 5784 3713 5818
rect 3747 5784 3781 5818
rect 3815 5784 3849 5818
rect 3883 5784 3917 5818
rect 3951 5784 3985 5818
rect 4019 5784 4053 5818
rect 4087 5784 4121 5818
rect 4155 5784 4189 5818
rect 4223 5784 4257 5818
rect 4291 5784 4325 5818
rect 4359 5784 4393 5818
rect 4427 5784 4461 5818
rect 4495 5784 4529 5818
rect 4563 5784 4597 5818
rect 4631 5784 4665 5818
rect 4699 5784 4733 5818
rect 4767 5784 4801 5818
rect 4835 5784 4869 5818
rect 4903 5784 4937 5818
rect 4971 5784 5005 5818
rect 5039 5784 5073 5818
rect 5107 5804 6781 5818
rect 5107 5798 6040 5804
rect 5107 5784 5155 5798
rect 3340 5764 5155 5784
rect 5189 5764 5223 5798
rect 5257 5764 5291 5798
rect 5325 5764 5359 5798
rect 5393 5764 5427 5798
rect 5461 5764 5495 5798
rect 5529 5764 5563 5798
rect 5597 5764 5631 5798
rect 5665 5764 5699 5798
rect 5733 5764 5767 5798
rect 5801 5764 5835 5798
rect 5869 5764 5903 5798
rect 5937 5764 5971 5798
rect 6005 5770 6040 5798
rect 6074 5770 6108 5804
rect 6142 5770 6176 5804
rect 6210 5770 6244 5804
rect 6278 5770 6312 5804
rect 6346 5770 6380 5804
rect 6414 5770 6448 5804
rect 6482 5770 6516 5804
rect 6550 5770 6584 5804
rect 6618 5770 6652 5804
rect 6686 5770 6720 5804
rect 6754 5770 6781 5804
rect 6005 5764 6781 5770
rect 3340 5748 6781 5764
rect 3340 5714 3373 5748
rect 3407 5714 3441 5748
rect 3475 5714 3509 5748
rect 3543 5714 3577 5748
rect 3611 5714 3645 5748
rect 3679 5714 3713 5748
rect 3747 5714 3781 5748
rect 3815 5714 3849 5748
rect 3883 5714 3917 5748
rect 3951 5714 3985 5748
rect 4019 5714 4053 5748
rect 4087 5714 4121 5748
rect 4155 5714 4189 5748
rect 4223 5714 4257 5748
rect 4291 5714 4325 5748
rect 4359 5714 4393 5748
rect 4427 5714 4461 5748
rect 4495 5714 4529 5748
rect 4563 5714 4597 5748
rect 4631 5714 4665 5748
rect 4699 5714 4733 5748
rect 4767 5714 4801 5748
rect 4835 5714 4869 5748
rect 4903 5714 4937 5748
rect 4971 5714 5005 5748
rect 5039 5714 5073 5748
rect 5107 5735 6781 5748
rect 5107 5728 6040 5735
rect 5107 5714 5155 5728
rect 3340 5694 5155 5714
rect 5189 5694 5223 5728
rect 5257 5694 5291 5728
rect 5325 5694 5359 5728
rect 5393 5694 5427 5728
rect 5461 5694 5495 5728
rect 5529 5694 5563 5728
rect 5597 5694 5631 5728
rect 5665 5694 5699 5728
rect 5733 5694 5767 5728
rect 5801 5694 5835 5728
rect 5869 5694 5903 5728
rect 5937 5694 5971 5728
rect 6005 5701 6040 5728
rect 6074 5701 6108 5735
rect 6142 5701 6176 5735
rect 6210 5701 6244 5735
rect 6278 5701 6312 5735
rect 6346 5701 6380 5735
rect 6414 5701 6448 5735
rect 6482 5701 6516 5735
rect 6550 5701 6584 5735
rect 6618 5701 6652 5735
rect 6686 5701 6720 5735
rect 6754 5723 6781 5735
rect 6754 5701 6825 5723
rect 6005 5694 6825 5701
rect 3340 5689 6825 5694
rect 6859 5689 6893 5723
rect 6927 5689 6961 5723
rect 6995 5689 7029 5723
rect 7063 5689 7097 5723
rect 7131 5689 7165 5723
rect 7199 5689 7233 5723
rect 7267 5689 7301 5723
rect 7335 5689 7369 5723
rect 7403 5689 7437 5723
rect 7471 5689 7505 5723
rect 7539 5689 7573 5723
rect 7607 5689 7641 5723
rect 7675 5689 7709 5723
rect 7743 5689 7777 5723
rect 7811 5689 7845 5723
rect 7879 5689 7913 5723
rect 7947 5689 7981 5723
rect 8015 5689 8049 5723
rect 8083 5689 8117 5723
rect 8151 5689 8185 5723
rect 8219 5689 8253 5723
rect 8287 5689 8321 5723
rect 8355 5689 8389 5723
rect 8423 5689 8457 5723
rect 8491 5689 8525 5723
rect 8559 5689 8593 5723
rect 8627 5689 8661 5723
rect 8695 5689 8729 5723
rect 8763 5689 8797 5723
rect 8831 5689 8865 5723
rect 8899 5689 8933 5723
rect 8967 5689 9001 5723
rect 9035 5689 9069 5723
rect 9103 5689 9137 5723
rect 9171 5689 9205 5723
rect 9239 5689 9273 5723
rect 9307 5689 9341 5723
rect 9375 5689 9409 5723
rect 9443 5689 9477 5723
rect 9511 5689 9545 5723
rect 9579 5689 9613 5723
rect 9647 5689 9681 5723
rect 9715 5689 9749 5723
rect 9783 5689 9817 5723
rect 9851 5689 9886 5723
rect 9920 5689 9955 5723
rect 9989 5689 10024 5723
rect 10058 5689 10093 5723
rect 10127 5689 10162 5723
rect 10196 5689 10231 5723
rect 10265 5689 10300 5723
rect 10334 5689 10369 5723
rect 10403 5689 10438 5723
rect 10472 5689 10507 5723
rect 10541 5689 10576 5723
rect 10610 5689 10645 5723
rect 10679 5689 10714 5723
rect 10748 5689 10783 5723
rect 10817 5689 10852 5723
rect 10886 5689 10921 5723
rect 10955 5689 10990 5723
rect 11024 5689 11059 5723
rect 11093 5689 11128 5723
rect 11162 5689 11197 5723
rect 11231 5689 11266 5723
rect 11300 5689 11335 5723
rect 11369 5689 11404 5723
rect 11438 5689 11473 5723
rect 11507 5689 11542 5723
rect 11576 5689 11611 5723
rect 11645 5689 11680 5723
rect 11714 5689 11749 5723
rect 11783 5689 11818 5723
rect 11852 5689 11887 5723
rect 11921 5689 11956 5723
rect 11990 5689 12025 5723
rect 12059 5689 12094 5723
rect 12128 5689 12163 5723
rect 12197 5689 12232 5723
rect 12266 5689 12301 5723
rect 12335 5689 12370 5723
rect 12404 5689 12439 5723
rect 12473 5689 12508 5723
rect 12542 5689 12577 5723
rect 12611 5689 12646 5723
rect 12680 5689 12715 5723
rect 12749 5689 12784 5723
rect 12818 5689 12853 5723
rect 12887 5689 12922 5723
rect 12956 5689 12991 5723
rect 13025 5689 13060 5723
rect 13094 5689 13129 5723
rect 13163 5689 13197 5723
rect 3340 5678 6781 5689
rect 3340 5644 3373 5678
rect 3407 5644 3441 5678
rect 3475 5644 3509 5678
rect 3543 5644 3577 5678
rect 3611 5644 3645 5678
rect 3679 5644 3713 5678
rect 3747 5644 3781 5678
rect 3815 5644 3849 5678
rect 3883 5644 3917 5678
rect 3951 5644 3985 5678
rect 4019 5644 4053 5678
rect 4087 5644 4121 5678
rect 4155 5644 4189 5678
rect 4223 5644 4257 5678
rect 4291 5644 4325 5678
rect 4359 5644 4393 5678
rect 4427 5644 4461 5678
rect 4495 5644 4529 5678
rect 4563 5644 4597 5678
rect 4631 5644 4665 5678
rect 4699 5644 4733 5678
rect 4767 5644 4801 5678
rect 4835 5644 4869 5678
rect 4903 5644 4937 5678
rect 4971 5644 5005 5678
rect 5039 5644 5073 5678
rect 5107 5666 6781 5678
rect 5107 5657 6040 5666
rect 5107 5644 5155 5657
rect 3340 5623 5155 5644
rect 5189 5623 5223 5657
rect 5257 5623 5291 5657
rect 5325 5623 5359 5657
rect 5393 5623 5427 5657
rect 5461 5623 5495 5657
rect 5529 5623 5563 5657
rect 5597 5623 5631 5657
rect 5665 5623 5699 5657
rect 5733 5623 5767 5657
rect 5801 5623 5835 5657
rect 5869 5623 5903 5657
rect 5937 5623 5971 5657
rect 6005 5632 6040 5657
rect 6074 5632 6108 5666
rect 6142 5632 6176 5666
rect 6210 5632 6244 5666
rect 6278 5632 6312 5666
rect 6346 5632 6380 5666
rect 6414 5632 6448 5666
rect 6482 5632 6516 5666
rect 6550 5632 6584 5666
rect 6618 5632 6652 5666
rect 6686 5632 6720 5666
rect 6754 5632 6781 5666
rect 6005 5623 6781 5632
rect 3340 5608 6781 5623
rect 3340 5574 3373 5608
rect 3407 5574 3441 5608
rect 3475 5574 3509 5608
rect 3543 5574 3577 5608
rect 3611 5574 3645 5608
rect 3679 5574 3713 5608
rect 3747 5574 3781 5608
rect 3815 5574 3849 5608
rect 3883 5574 3917 5608
rect 3951 5574 3985 5608
rect 4019 5574 4053 5608
rect 4087 5574 4121 5608
rect 4155 5574 4189 5608
rect 4223 5574 4257 5608
rect 4291 5574 4325 5608
rect 4359 5574 4393 5608
rect 4427 5574 4461 5608
rect 4495 5574 4529 5608
rect 4563 5574 4597 5608
rect 4631 5574 4665 5608
rect 4699 5574 4733 5608
rect 4767 5574 4801 5608
rect 4835 5574 4869 5608
rect 4903 5574 4937 5608
rect 4971 5574 5005 5608
rect 5039 5574 5073 5608
rect 5107 5597 6781 5608
rect 5107 5586 6040 5597
rect 5107 5574 5155 5586
rect 3340 5552 5155 5574
rect 5189 5552 5223 5586
rect 5257 5552 5291 5586
rect 5325 5552 5359 5586
rect 5393 5552 5427 5586
rect 5461 5552 5495 5586
rect 5529 5552 5563 5586
rect 5597 5552 5631 5586
rect 5665 5552 5699 5586
rect 5733 5552 5767 5586
rect 5801 5552 5835 5586
rect 5869 5552 5903 5586
rect 5937 5552 5971 5586
rect 6005 5563 6040 5586
rect 6074 5563 6108 5597
rect 6142 5563 6176 5597
rect 6210 5563 6244 5597
rect 6278 5563 6312 5597
rect 6346 5563 6380 5597
rect 6414 5563 6448 5597
rect 6482 5563 6516 5597
rect 6550 5563 6584 5597
rect 6618 5563 6652 5597
rect 6686 5563 6720 5597
rect 6754 5563 6781 5597
rect 6005 5552 6781 5563
rect 3340 5538 6781 5552
rect 3340 5504 3373 5538
rect 3407 5504 3441 5538
rect 3475 5504 3509 5538
rect 3543 5504 3577 5538
rect 3611 5504 3645 5538
rect 3679 5504 3713 5538
rect 3747 5504 3781 5538
rect 3815 5504 3849 5538
rect 3883 5504 3917 5538
rect 3951 5504 3985 5538
rect 4019 5504 4053 5538
rect 4087 5504 4121 5538
rect 4155 5504 4189 5538
rect 4223 5504 4257 5538
rect 4291 5504 4325 5538
rect 4359 5504 4393 5538
rect 4427 5504 4461 5538
rect 4495 5504 4529 5538
rect 4563 5504 4597 5538
rect 4631 5504 4665 5538
rect 4699 5504 4733 5538
rect 4767 5504 4801 5538
rect 4835 5504 4869 5538
rect 4903 5504 4937 5538
rect 4971 5504 5005 5538
rect 5039 5504 5073 5538
rect 5107 5528 6781 5538
rect 5107 5505 6040 5528
rect 5107 5504 5155 5505
rect 3340 5471 5155 5504
rect 5189 5471 5223 5505
rect 5257 5471 5291 5505
rect 5325 5471 5359 5505
rect 5393 5471 5427 5505
rect 5461 5471 5495 5505
rect 5529 5471 5563 5505
rect 5597 5471 5631 5505
rect 5665 5471 5699 5505
rect 5733 5471 5767 5505
rect 5801 5471 5835 5505
rect 5869 5471 5903 5505
rect 5937 5471 5971 5505
rect 6005 5494 6040 5505
rect 6074 5494 6108 5528
rect 6142 5494 6176 5528
rect 6210 5494 6244 5528
rect 6278 5494 6312 5528
rect 6346 5494 6380 5528
rect 6414 5494 6448 5528
rect 6482 5494 6516 5528
rect 6550 5494 6584 5528
rect 6618 5494 6652 5528
rect 6686 5494 6720 5528
rect 6754 5494 6781 5528
rect 6005 5471 6781 5494
rect 3340 5468 6781 5471
rect 3340 5434 3373 5468
rect 3407 5434 3441 5468
rect 3475 5434 3509 5468
rect 3543 5434 3577 5468
rect 3611 5434 3645 5468
rect 3679 5434 3713 5468
rect 3747 5434 3781 5468
rect 3815 5434 3849 5468
rect 3883 5434 3917 5468
rect 3951 5434 3985 5468
rect 4019 5434 4053 5468
rect 4087 5434 4121 5468
rect 4155 5434 4189 5468
rect 4223 5434 4257 5468
rect 4291 5434 4325 5468
rect 4359 5434 4393 5468
rect 4427 5434 4461 5468
rect 4495 5434 4529 5468
rect 4563 5434 4597 5468
rect 4631 5434 4665 5468
rect 4699 5434 4733 5468
rect 4767 5434 4801 5468
rect 4835 5434 4869 5468
rect 4903 5434 4937 5468
rect 4971 5434 5005 5468
rect 5039 5434 5073 5468
rect 5107 5459 6781 5468
rect 5107 5434 6040 5459
rect 3340 5431 6040 5434
rect 3340 5398 5155 5431
rect 3340 5364 3373 5398
rect 3407 5364 3441 5398
rect 3475 5364 3509 5398
rect 3543 5364 3577 5398
rect 3611 5364 3645 5398
rect 3679 5364 3713 5398
rect 3747 5364 3781 5398
rect 3815 5364 3849 5398
rect 3883 5364 3917 5398
rect 3951 5364 3985 5398
rect 4019 5364 4053 5398
rect 4087 5364 4121 5398
rect 4155 5364 4189 5398
rect 4223 5364 4257 5398
rect 4291 5364 4325 5398
rect 4359 5364 4393 5398
rect 4427 5364 4461 5398
rect 4495 5364 4529 5398
rect 4563 5364 4597 5398
rect 4631 5364 4665 5398
rect 4699 5364 4733 5398
rect 4767 5364 4801 5398
rect 4835 5364 4869 5398
rect 4903 5364 4937 5398
rect 4971 5364 5005 5398
rect 5039 5364 5073 5398
rect 5107 5397 5155 5398
rect 5189 5397 5223 5431
rect 5257 5397 5291 5431
rect 5325 5397 5359 5431
rect 5393 5397 5427 5431
rect 5461 5397 5495 5431
rect 5529 5397 5563 5431
rect 5597 5397 5631 5431
rect 5665 5397 5699 5431
rect 5733 5397 5767 5431
rect 5801 5397 5835 5431
rect 5869 5397 5903 5431
rect 5937 5397 5971 5431
rect 6005 5425 6040 5431
rect 6074 5425 6108 5459
rect 6142 5425 6176 5459
rect 6210 5425 6244 5459
rect 6278 5425 6312 5459
rect 6346 5425 6380 5459
rect 6414 5425 6448 5459
rect 6482 5425 6516 5459
rect 6550 5425 6584 5459
rect 6618 5425 6652 5459
rect 6686 5425 6720 5459
rect 6754 5425 6781 5459
rect 6005 5397 6781 5425
rect 5107 5390 6781 5397
rect 5107 5364 6040 5390
rect 3340 5356 6040 5364
rect 6074 5356 6108 5390
rect 6142 5356 6176 5390
rect 6210 5356 6244 5390
rect 6278 5356 6312 5390
rect 6346 5356 6380 5390
rect 6414 5356 6448 5390
rect 6482 5356 6516 5390
rect 6550 5356 6584 5390
rect 6618 5356 6652 5390
rect 6686 5356 6720 5390
rect 6754 5375 6781 5390
rect 6754 5356 6825 5375
rect 3340 5328 5155 5356
rect 3340 5294 3373 5328
rect 3407 5294 3441 5328
rect 3475 5294 3509 5328
rect 3543 5294 3577 5328
rect 3611 5294 3645 5328
rect 3679 5294 3713 5328
rect 3747 5294 3781 5328
rect 3815 5294 3849 5328
rect 3883 5294 3917 5328
rect 3951 5294 3985 5328
rect 4019 5294 4053 5328
rect 4087 5294 4121 5328
rect 4155 5294 4189 5328
rect 4223 5294 4257 5328
rect 4291 5294 4325 5328
rect 4359 5294 4393 5328
rect 4427 5294 4461 5328
rect 4495 5294 4529 5328
rect 4563 5294 4597 5328
rect 4631 5294 4665 5328
rect 4699 5294 4733 5328
rect 4767 5294 4801 5328
rect 4835 5294 4869 5328
rect 4903 5294 4937 5328
rect 4971 5294 5005 5328
rect 5039 5294 5073 5328
rect 5107 5322 5155 5328
rect 5189 5322 5223 5356
rect 5257 5322 5291 5356
rect 5325 5322 5359 5356
rect 5393 5322 5427 5356
rect 5461 5322 5495 5356
rect 5529 5322 5563 5356
rect 5597 5322 5631 5356
rect 5665 5322 5699 5356
rect 5733 5322 5767 5356
rect 5801 5322 5835 5356
rect 5869 5322 5903 5356
rect 5937 5322 5971 5356
rect 6005 5341 6825 5356
rect 6859 5341 6893 5375
rect 6927 5341 6961 5375
rect 6995 5341 7029 5375
rect 7063 5341 7097 5375
rect 7131 5341 7165 5375
rect 7199 5341 7233 5375
rect 7267 5341 7301 5375
rect 7335 5341 7369 5375
rect 7403 5341 7437 5375
rect 7471 5341 7505 5375
rect 7539 5341 7573 5375
rect 7607 5341 7641 5375
rect 7675 5341 7709 5375
rect 7743 5341 7777 5375
rect 7811 5341 7845 5375
rect 7879 5341 7913 5375
rect 7947 5341 7981 5375
rect 8015 5341 8049 5375
rect 8083 5341 8117 5375
rect 8151 5341 8185 5375
rect 8219 5341 8253 5375
rect 8287 5341 8321 5375
rect 8355 5341 8389 5375
rect 8423 5341 8457 5375
rect 8491 5341 8525 5375
rect 8559 5341 8593 5375
rect 8627 5341 8661 5375
rect 8695 5341 8729 5375
rect 8763 5341 8797 5375
rect 8831 5341 8865 5375
rect 8899 5341 8933 5375
rect 8967 5341 9001 5375
rect 9035 5341 9069 5375
rect 9103 5341 9137 5375
rect 9171 5341 9205 5375
rect 9239 5341 9273 5375
rect 9307 5341 9341 5375
rect 9375 5341 9409 5375
rect 9443 5341 9477 5375
rect 9511 5341 9545 5375
rect 9579 5341 9613 5375
rect 9647 5341 9681 5375
rect 9715 5341 9749 5375
rect 9783 5341 9817 5375
rect 9851 5341 9886 5375
rect 9920 5341 9955 5375
rect 9989 5341 10024 5375
rect 10058 5341 10093 5375
rect 10127 5341 10162 5375
rect 10196 5341 10231 5375
rect 10265 5341 10300 5375
rect 10334 5341 10369 5375
rect 10403 5341 10438 5375
rect 10472 5341 10507 5375
rect 10541 5341 10576 5375
rect 10610 5341 10645 5375
rect 10679 5341 10714 5375
rect 10748 5341 10783 5375
rect 10817 5341 10852 5375
rect 10886 5341 10921 5375
rect 10955 5341 10990 5375
rect 11024 5341 11059 5375
rect 11093 5341 11128 5375
rect 11162 5341 11197 5375
rect 11231 5341 11266 5375
rect 11300 5341 11335 5375
rect 11369 5341 11404 5375
rect 11438 5341 11473 5375
rect 11507 5341 11542 5375
rect 11576 5341 11611 5375
rect 11645 5341 11680 5375
rect 11714 5341 11749 5375
rect 11783 5341 11818 5375
rect 11852 5341 11887 5375
rect 11921 5341 11956 5375
rect 11990 5341 12025 5375
rect 12059 5341 12094 5375
rect 12128 5341 12163 5375
rect 12197 5341 12232 5375
rect 12266 5341 12301 5375
rect 12335 5341 12370 5375
rect 12404 5341 12439 5375
rect 12473 5341 12508 5375
rect 12542 5341 12577 5375
rect 12611 5341 12646 5375
rect 12680 5341 12715 5375
rect 12749 5341 12784 5375
rect 12818 5341 12853 5375
rect 12887 5341 12922 5375
rect 12956 5341 12991 5375
rect 13025 5341 13060 5375
rect 13094 5341 13129 5375
rect 13163 5341 13197 5375
rect 6005 5322 6781 5341
rect 5107 5321 6781 5322
rect 5107 5294 6040 5321
rect 3340 5287 6040 5294
rect 6074 5287 6108 5321
rect 6142 5287 6176 5321
rect 6210 5287 6244 5321
rect 6278 5287 6312 5321
rect 6346 5287 6380 5321
rect 6414 5287 6448 5321
rect 6482 5287 6516 5321
rect 6550 5287 6584 5321
rect 6618 5287 6652 5321
rect 6686 5287 6720 5321
rect 6754 5287 6781 5321
rect 3340 5281 6781 5287
rect 3340 5257 5155 5281
rect 3340 5223 3373 5257
rect 3407 5223 3441 5257
rect 3475 5223 3509 5257
rect 3543 5223 3577 5257
rect 3611 5223 3645 5257
rect 3679 5223 3713 5257
rect 3747 5223 3781 5257
rect 3815 5223 3849 5257
rect 3883 5223 3917 5257
rect 3951 5223 3985 5257
rect 4019 5223 4053 5257
rect 4087 5223 4121 5257
rect 4155 5223 4189 5257
rect 4223 5223 4257 5257
rect 4291 5223 4325 5257
rect 4359 5223 4393 5257
rect 4427 5223 4461 5257
rect 4495 5223 4529 5257
rect 4563 5223 4597 5257
rect 4631 5223 4665 5257
rect 4699 5223 4733 5257
rect 4767 5223 4801 5257
rect 4835 5223 4869 5257
rect 4903 5223 4937 5257
rect 4971 5223 5005 5257
rect 5039 5223 5073 5257
rect 5107 5247 5155 5257
rect 5189 5247 5223 5281
rect 5257 5247 5291 5281
rect 5325 5247 5359 5281
rect 5393 5247 5427 5281
rect 5461 5247 5495 5281
rect 5529 5247 5563 5281
rect 5597 5247 5631 5281
rect 5665 5247 5699 5281
rect 5733 5247 5767 5281
rect 5801 5247 5835 5281
rect 5869 5247 5903 5281
rect 5937 5247 5971 5281
rect 6005 5251 6781 5281
rect 6005 5247 6040 5251
rect 5107 5223 6040 5247
rect 3340 5217 6040 5223
rect 6074 5217 6108 5251
rect 6142 5217 6176 5251
rect 6210 5217 6244 5251
rect 6278 5217 6312 5251
rect 6346 5217 6380 5251
rect 6414 5217 6448 5251
rect 6482 5217 6516 5251
rect 6550 5217 6584 5251
rect 6618 5217 6652 5251
rect 6686 5217 6720 5251
rect 6754 5217 6781 5251
rect 3340 5206 6781 5217
rect 3340 5186 5155 5206
rect 3340 5152 3373 5186
rect 3407 5152 3441 5186
rect 3475 5152 3509 5186
rect 3543 5152 3577 5186
rect 3611 5152 3645 5186
rect 3679 5152 3713 5186
rect 3747 5152 3781 5186
rect 3815 5152 3849 5186
rect 3883 5152 3917 5186
rect 3951 5152 3985 5186
rect 4019 5152 4053 5186
rect 4087 5152 4121 5186
rect 4155 5152 4189 5186
rect 4223 5152 4257 5186
rect 4291 5152 4325 5186
rect 4359 5152 4393 5186
rect 4427 5152 4461 5186
rect 4495 5152 4529 5186
rect 4563 5152 4597 5186
rect 4631 5152 4665 5186
rect 4699 5152 4733 5186
rect 4767 5152 4801 5186
rect 4835 5152 4869 5186
rect 4903 5152 4937 5186
rect 4971 5152 5005 5186
rect 5039 5152 5073 5186
rect 5107 5172 5155 5186
rect 5189 5172 5223 5206
rect 5257 5172 5291 5206
rect 5325 5172 5359 5206
rect 5393 5172 5427 5206
rect 5461 5172 5495 5206
rect 5529 5172 5563 5206
rect 5597 5172 5631 5206
rect 5665 5172 5699 5206
rect 5733 5172 5767 5206
rect 5801 5172 5835 5206
rect 5869 5172 5903 5206
rect 5937 5172 5971 5206
rect 6005 5181 6781 5206
rect 6005 5172 6040 5181
rect 5107 5152 6040 5172
rect 3340 5147 6040 5152
rect 6074 5147 6108 5181
rect 6142 5147 6176 5181
rect 6210 5147 6244 5181
rect 6278 5147 6312 5181
rect 6346 5147 6380 5181
rect 6414 5147 6448 5181
rect 6482 5147 6516 5181
rect 6550 5147 6584 5181
rect 6618 5147 6652 5181
rect 6686 5147 6720 5181
rect 6754 5147 6781 5181
rect 3340 5131 6781 5147
rect 3340 5115 5155 5131
rect 3340 5081 3373 5115
rect 3407 5081 3441 5115
rect 3475 5081 3509 5115
rect 3543 5081 3577 5115
rect 3611 5081 3645 5115
rect 3679 5081 3713 5115
rect 3747 5081 3781 5115
rect 3815 5081 3849 5115
rect 3883 5081 3917 5115
rect 3951 5081 3985 5115
rect 4019 5081 4053 5115
rect 4087 5081 4121 5115
rect 4155 5081 4189 5115
rect 4223 5081 4257 5115
rect 4291 5081 4325 5115
rect 4359 5081 4393 5115
rect 4427 5081 4461 5115
rect 4495 5081 4529 5115
rect 4563 5081 4597 5115
rect 4631 5081 4665 5115
rect 4699 5081 4733 5115
rect 4767 5081 4801 5115
rect 4835 5081 4869 5115
rect 4903 5081 4937 5115
rect 4971 5081 5005 5115
rect 5039 5081 5073 5115
rect 5107 5097 5155 5115
rect 5189 5097 5223 5131
rect 5257 5097 5291 5131
rect 5325 5097 5359 5131
rect 5393 5097 5427 5131
rect 5461 5097 5495 5131
rect 5529 5097 5563 5131
rect 5597 5097 5631 5131
rect 5665 5097 5699 5131
rect 5733 5097 5767 5131
rect 5801 5097 5835 5131
rect 5869 5097 5903 5131
rect 5937 5097 5971 5131
rect 6005 5111 6781 5131
rect 6005 5097 6040 5111
rect 5107 5081 6040 5097
rect 3340 5077 6040 5081
rect 6074 5077 6108 5111
rect 6142 5077 6176 5111
rect 6210 5077 6244 5111
rect 6278 5077 6312 5111
rect 6346 5077 6380 5111
rect 6414 5077 6448 5111
rect 6482 5077 6516 5111
rect 6550 5077 6584 5111
rect 6618 5077 6652 5111
rect 6686 5077 6720 5111
rect 6754 5077 6781 5111
rect 3340 5056 6781 5077
rect 3340 5044 5155 5056
rect 3340 5010 3373 5044
rect 3407 5010 3441 5044
rect 3475 5010 3509 5044
rect 3543 5010 3577 5044
rect 3611 5010 3645 5044
rect 3679 5010 3713 5044
rect 3747 5010 3781 5044
rect 3815 5010 3849 5044
rect 3883 5010 3917 5044
rect 3951 5010 3985 5044
rect 4019 5010 4053 5044
rect 4087 5010 4121 5044
rect 4155 5010 4189 5044
rect 4223 5010 4257 5044
rect 4291 5010 4325 5044
rect 4359 5010 4393 5044
rect 4427 5010 4461 5044
rect 4495 5010 4529 5044
rect 4563 5010 4597 5044
rect 4631 5010 4665 5044
rect 4699 5010 4733 5044
rect 4767 5010 4801 5044
rect 4835 5010 4869 5044
rect 4903 5010 4937 5044
rect 4971 5010 5005 5044
rect 5039 5010 5073 5044
rect 5107 5022 5155 5044
rect 5189 5022 5223 5056
rect 5257 5022 5291 5056
rect 5325 5022 5359 5056
rect 5393 5022 5427 5056
rect 5461 5022 5495 5056
rect 5529 5022 5563 5056
rect 5597 5022 5631 5056
rect 5665 5022 5699 5056
rect 5733 5022 5767 5056
rect 5801 5022 5835 5056
rect 5869 5022 5903 5056
rect 5937 5022 5971 5056
rect 6005 5041 6781 5056
rect 6005 5022 6040 5041
rect 5107 5010 6040 5022
rect 3340 5007 6040 5010
rect 6074 5007 6108 5041
rect 6142 5007 6176 5041
rect 6210 5007 6244 5041
rect 6278 5007 6312 5041
rect 6346 5007 6380 5041
rect 6414 5007 6448 5041
rect 6482 5007 6516 5041
rect 6550 5007 6584 5041
rect 6618 5007 6652 5041
rect 6686 5007 6720 5041
rect 6754 5007 6781 5041
rect 3340 4985 6781 5007
rect 3340 4981 6829 4985
rect 3340 4973 5155 4981
rect 3340 4939 3373 4973
rect 3407 4939 3441 4973
rect 3475 4939 3509 4973
rect 3543 4939 3577 4973
rect 3611 4939 3645 4973
rect 3679 4939 3713 4973
rect 3747 4939 3781 4973
rect 3815 4939 3849 4973
rect 3883 4939 3917 4973
rect 3951 4939 3985 4973
rect 4019 4939 4053 4973
rect 4087 4939 4121 4973
rect 4155 4939 4189 4973
rect 4223 4939 4257 4973
rect 4291 4939 4325 4973
rect 4359 4939 4393 4973
rect 4427 4939 4461 4973
rect 4495 4939 4529 4973
rect 4563 4939 4597 4973
rect 4631 4939 4665 4973
rect 4699 4939 4733 4973
rect 4767 4939 4801 4973
rect 4835 4939 4869 4973
rect 4903 4939 4937 4973
rect 4971 4939 5005 4973
rect 5039 4939 5073 4973
rect 5107 4947 5155 4973
rect 5189 4947 5223 4981
rect 5257 4947 5291 4981
rect 5325 4947 5359 4981
rect 5393 4947 5427 4981
rect 5461 4947 5495 4981
rect 5529 4947 5563 4981
rect 5597 4947 5631 4981
rect 5665 4947 5699 4981
rect 5733 4947 5767 4981
rect 5801 4947 5835 4981
rect 5869 4947 5903 4981
rect 5937 4947 5971 4981
rect 6005 4971 6829 4981
rect 6005 4947 6040 4971
rect 5107 4939 6040 4947
rect 3340 4937 6040 4939
rect 6074 4937 6108 4971
rect 6142 4937 6176 4971
rect 6210 4937 6244 4971
rect 6278 4937 6312 4971
rect 6346 4937 6380 4971
rect 6414 4937 6448 4971
rect 6482 4937 6516 4971
rect 6550 4937 6584 4971
rect 6618 4937 6652 4971
rect 6686 4937 6720 4971
rect 6754 4951 6829 4971
rect 6863 4951 6898 4985
rect 6932 4951 6967 4985
rect 7001 4951 7036 4985
rect 7070 4951 7105 4985
rect 7139 4951 7174 4985
rect 7208 4951 7243 4985
rect 7277 4951 7312 4985
rect 7346 4951 7381 4985
rect 7415 4951 7450 4985
rect 7484 4951 7519 4985
rect 7553 4951 7588 4985
rect 7622 4951 7657 4985
rect 7691 4951 7726 4985
rect 7760 4951 7795 4985
rect 7829 4951 7864 4985
rect 7898 4951 7933 4985
rect 7967 4951 8002 4985
rect 8036 4951 8071 4985
rect 8105 4951 8140 4985
rect 8174 4951 8209 4985
rect 8243 4951 8278 4985
rect 8312 4951 8347 4985
rect 8381 4951 8416 4985
rect 8450 4951 8485 4985
rect 8519 4951 8554 4985
rect 8588 4951 8623 4985
rect 6754 4937 8623 4951
rect 3340 4917 8623 4937
rect 3340 4906 6829 4917
rect 3340 4902 5155 4906
rect 3340 4868 3373 4902
rect 3407 4868 3441 4902
rect 3475 4868 3509 4902
rect 3543 4868 3577 4902
rect 3611 4868 3645 4902
rect 3679 4868 3713 4902
rect 3747 4868 3781 4902
rect 3815 4868 3849 4902
rect 3883 4868 3917 4902
rect 3951 4868 3985 4902
rect 4019 4868 4053 4902
rect 4087 4868 4121 4902
rect 4155 4868 4189 4902
rect 4223 4868 4257 4902
rect 4291 4868 4325 4902
rect 4359 4868 4393 4902
rect 4427 4868 4461 4902
rect 4495 4868 4529 4902
rect 4563 4868 4597 4902
rect 4631 4868 4665 4902
rect 4699 4868 4733 4902
rect 4767 4868 4801 4902
rect 4835 4868 4869 4902
rect 4903 4868 4937 4902
rect 4971 4868 5005 4902
rect 5039 4868 5073 4902
rect 5107 4872 5155 4902
rect 5189 4872 5223 4906
rect 5257 4872 5291 4906
rect 5325 4872 5359 4906
rect 5393 4872 5427 4906
rect 5461 4872 5495 4906
rect 5529 4872 5563 4906
rect 5597 4872 5631 4906
rect 5665 4872 5699 4906
rect 5733 4872 5767 4906
rect 5801 4872 5835 4906
rect 5869 4872 5903 4906
rect 5937 4872 5971 4906
rect 6005 4901 6829 4906
rect 6005 4872 6040 4901
rect 5107 4868 6040 4872
rect 3340 4867 6040 4868
rect 6074 4867 6108 4901
rect 6142 4867 6176 4901
rect 6210 4867 6244 4901
rect 6278 4867 6312 4901
rect 6346 4867 6380 4901
rect 6414 4867 6448 4901
rect 6482 4867 6516 4901
rect 6550 4867 6584 4901
rect 6618 4867 6652 4901
rect 6686 4867 6720 4901
rect 6754 4883 6829 4901
rect 6863 4883 6898 4917
rect 6932 4883 6967 4917
rect 7001 4883 7036 4917
rect 7070 4883 7105 4917
rect 7139 4883 7174 4917
rect 7208 4883 7243 4917
rect 7277 4883 7312 4917
rect 7346 4883 7381 4917
rect 7415 4883 7450 4917
rect 7484 4883 7519 4917
rect 7553 4883 7588 4917
rect 7622 4883 7657 4917
rect 7691 4883 7726 4917
rect 7760 4883 7795 4917
rect 7829 4883 7864 4917
rect 7898 4883 7933 4917
rect 7967 4883 8002 4917
rect 8036 4883 8071 4917
rect 8105 4883 8140 4917
rect 8174 4883 8209 4917
rect 8243 4883 8278 4917
rect 8312 4883 8347 4917
rect 8381 4883 8416 4917
rect 8450 4883 8485 4917
rect 8519 4883 8554 4917
rect 8588 4883 8623 4917
rect 6754 4867 8623 4883
rect 3340 4849 8623 4867
rect 3340 4831 6829 4849
rect 3340 4797 3373 4831
rect 3407 4797 3441 4831
rect 3475 4797 3509 4831
rect 3543 4797 3577 4831
rect 3611 4797 3645 4831
rect 3679 4797 3713 4831
rect 3747 4797 3781 4831
rect 3815 4797 3849 4831
rect 3883 4797 3917 4831
rect 3951 4797 3985 4831
rect 4019 4797 4053 4831
rect 4087 4797 4121 4831
rect 4155 4797 4189 4831
rect 4223 4797 4257 4831
rect 4291 4797 4325 4831
rect 4359 4797 4393 4831
rect 4427 4797 4461 4831
rect 4495 4797 4529 4831
rect 4563 4797 4597 4831
rect 4631 4797 4665 4831
rect 4699 4797 4733 4831
rect 4767 4797 4801 4831
rect 4835 4797 4869 4831
rect 4903 4797 4937 4831
rect 4971 4797 5005 4831
rect 5039 4797 5073 4831
rect 5107 4797 5155 4831
rect 5189 4797 5223 4831
rect 5257 4797 5291 4831
rect 5325 4797 5359 4831
rect 5393 4797 5427 4831
rect 5461 4797 5495 4831
rect 5529 4797 5563 4831
rect 5597 4797 5631 4831
rect 5665 4797 5699 4831
rect 5733 4797 5767 4831
rect 5801 4797 5835 4831
rect 5869 4797 5903 4831
rect 5937 4797 5971 4831
rect 6005 4797 6040 4831
rect 6074 4797 6108 4831
rect 6142 4797 6176 4831
rect 6210 4797 6244 4831
rect 6278 4797 6312 4831
rect 6346 4797 6380 4831
rect 6414 4797 6448 4831
rect 6482 4797 6516 4831
rect 6550 4797 6584 4831
rect 6618 4797 6652 4831
rect 6686 4797 6720 4831
rect 6754 4815 6829 4831
rect 6863 4815 6898 4849
rect 6932 4815 6967 4849
rect 7001 4815 7036 4849
rect 7070 4815 7105 4849
rect 7139 4815 7174 4849
rect 7208 4815 7243 4849
rect 7277 4815 7312 4849
rect 7346 4815 7381 4849
rect 7415 4815 7450 4849
rect 7484 4815 7519 4849
rect 7553 4815 7588 4849
rect 7622 4815 7657 4849
rect 7691 4815 7726 4849
rect 7760 4815 7795 4849
rect 7829 4815 7864 4849
rect 7898 4815 7933 4849
rect 7967 4815 8002 4849
rect 8036 4815 8071 4849
rect 8105 4815 8140 4849
rect 8174 4815 8209 4849
rect 8243 4815 8278 4849
rect 8312 4815 8347 4849
rect 8381 4815 8416 4849
rect 8450 4815 8485 4849
rect 8519 4815 8554 4849
rect 8588 4815 8623 4849
rect 13145 4815 13197 4985
rect 6754 4798 13197 4815
rect 6754 4797 13265 4798
rect 3340 4763 13265 4797
rect 3340 4729 3374 4763
rect 3408 4729 3443 4763
rect 3477 4729 3512 4763
rect 3546 4729 3581 4763
rect 3615 4729 3650 4763
rect 3684 4729 3719 4763
rect 3753 4729 3788 4763
rect 3822 4729 3857 4763
rect 3891 4729 3926 4763
rect 3960 4729 3995 4763
rect 4029 4729 4064 4763
rect 4098 4729 4133 4763
rect 4167 4729 4202 4763
rect 4236 4729 4271 4763
rect 4305 4729 4340 4763
rect 4374 4729 4409 4763
rect 4443 4729 4478 4763
rect 4512 4729 4547 4763
rect 4581 4729 4616 4763
rect 4650 4729 4685 4763
rect 4719 4729 4754 4763
rect 4788 4729 4823 4763
rect 4857 4729 4892 4763
rect 4926 4729 4961 4763
rect 4995 4729 5030 4763
rect 5064 4729 5099 4763
rect 5133 4729 5168 4763
rect 5202 4729 5237 4763
rect 5271 4729 5306 4763
rect 5340 4729 5375 4763
rect 5409 4729 5444 4763
rect 5478 4729 5513 4763
rect 5547 4729 5582 4763
rect 5616 4729 5651 4763
rect 5685 4729 5720 4763
rect 5754 4729 5789 4763
rect 5823 4729 5858 4763
rect 5892 4729 5927 4763
rect 5961 4729 5996 4763
rect 6030 4729 6065 4763
rect 6099 4729 6134 4763
rect 6168 4729 6203 4763
rect 6237 4729 6272 4763
rect 6306 4729 6341 4763
rect 6375 4729 6410 4763
rect 6444 4729 6479 4763
rect 6513 4729 6548 4763
rect 6582 4729 6617 4763
rect 6651 4729 6686 4763
rect 6720 4729 6755 4763
rect 6789 4729 6824 4763
rect 6858 4729 6893 4763
rect 6927 4729 6962 4763
rect 3340 4695 6962 4729
rect 10056 4729 10092 4763
rect 10126 4729 10161 4763
rect 10195 4729 10230 4763
rect 10264 4729 10299 4763
rect 10333 4729 10368 4763
rect 10402 4729 10437 4763
rect 10471 4729 10506 4763
rect 10540 4729 10575 4763
rect 10609 4729 10644 4763
rect 10678 4729 10713 4763
rect 10747 4729 10782 4763
rect 10816 4729 10851 4763
rect 10885 4729 10920 4763
rect 10954 4729 10989 4763
rect 11023 4729 11058 4763
rect 11092 4729 11127 4763
rect 11161 4729 11196 4763
rect 11230 4729 11265 4763
rect 11299 4729 11334 4763
rect 11368 4729 11403 4763
rect 11437 4729 11472 4763
rect 11506 4729 11541 4763
rect 11575 4729 11610 4763
rect 11644 4729 11679 4763
rect 11713 4729 11748 4763
rect 11782 4729 11817 4763
rect 11851 4729 11886 4763
rect 11920 4729 11955 4763
rect 11989 4729 12024 4763
rect 12058 4729 12093 4763
rect 12127 4729 12162 4763
rect 12196 4729 12231 4763
rect 12265 4729 12300 4763
rect 12334 4729 12369 4763
rect 12403 4729 12438 4763
rect 12472 4729 12507 4763
rect 12541 4729 12576 4763
rect 12610 4729 12645 4763
rect 12679 4729 12714 4763
rect 12748 4729 12783 4763
rect 12817 4729 12852 4763
rect 12886 4729 12921 4763
rect 12955 4729 12990 4763
rect 13024 4729 13059 4763
rect 13093 4729 13128 4763
rect 13162 4729 13197 4763
rect 13231 4730 13265 4763
rect 13231 4729 13333 4730
rect 10056 4696 13333 4729
rect 10056 4695 13367 4696
rect 3340 4661 3408 4695
rect 3442 4661 3477 4695
rect 3511 4661 3546 4695
rect 3580 4661 3615 4695
rect 3649 4661 3684 4695
rect 3718 4661 3753 4695
rect 3787 4661 3822 4695
rect 3856 4661 3891 4695
rect 3925 4661 3960 4695
rect 3994 4661 4029 4695
rect 4063 4661 4098 4695
rect 4132 4661 4167 4695
rect 4201 4661 4236 4695
rect 4270 4661 4305 4695
rect 4339 4661 4374 4695
rect 4408 4661 4443 4695
rect 4477 4661 4512 4695
rect 4546 4661 4581 4695
rect 4615 4661 4650 4695
rect 4684 4661 4718 4695
rect 3340 4657 4718 4661
rect 3374 4627 4718 4657
rect 3374 4623 3476 4627
rect 3340 4622 3476 4623
rect 3340 4588 3408 4622
rect 3442 4593 3476 4622
rect 3510 4593 3545 4627
rect 3579 4593 3614 4627
rect 3648 4593 3683 4627
rect 3717 4593 3752 4627
rect 3786 4593 3821 4627
rect 3855 4593 3890 4627
rect 3924 4593 3959 4627
rect 3993 4593 4028 4627
rect 4062 4593 4097 4627
rect 4131 4593 4166 4627
rect 4200 4593 4235 4627
rect 4269 4593 4304 4627
rect 4338 4593 4373 4627
rect 4407 4593 4442 4627
rect 4476 4593 4511 4627
rect 4545 4593 4580 4627
rect 4614 4593 4649 4627
rect 4683 4593 4718 4627
rect 10056 4661 10091 4695
rect 10125 4661 10160 4695
rect 10194 4661 10229 4695
rect 10263 4661 10298 4695
rect 10332 4661 10367 4695
rect 10401 4661 10436 4695
rect 10470 4661 10505 4695
rect 10539 4661 10574 4695
rect 10608 4661 10643 4695
rect 10677 4661 10712 4695
rect 10746 4661 10781 4695
rect 10815 4661 10850 4695
rect 10884 4661 10919 4695
rect 10953 4661 10988 4695
rect 11022 4661 11057 4695
rect 11091 4661 11126 4695
rect 11160 4661 11195 4695
rect 11229 4661 11264 4695
rect 11298 4661 11333 4695
rect 11367 4661 11402 4695
rect 11436 4661 11471 4695
rect 11505 4661 11540 4695
rect 11574 4661 11609 4695
rect 11643 4661 11678 4695
rect 11712 4661 11747 4695
rect 11781 4661 11816 4695
rect 11850 4661 11885 4695
rect 11919 4661 11954 4695
rect 11988 4661 12023 4695
rect 12057 4661 12092 4695
rect 12126 4661 12161 4695
rect 12195 4661 12230 4695
rect 12264 4661 12299 4695
rect 12333 4661 12368 4695
rect 12402 4661 12437 4695
rect 12471 4661 12506 4695
rect 12540 4661 12575 4695
rect 12609 4661 12644 4695
rect 12678 4661 12713 4695
rect 12747 4661 12782 4695
rect 12816 4661 12851 4695
rect 12885 4661 12920 4695
rect 12954 4661 12989 4695
rect 13023 4661 13058 4695
rect 13092 4661 13127 4695
rect 13161 4661 13196 4695
rect 13230 4661 13265 4695
rect 13299 4661 13367 4695
rect 10056 4627 13333 4661
rect 10056 4593 10091 4627
rect 10125 4593 10160 4627
rect 10194 4593 10229 4627
rect 10263 4593 10298 4627
rect 10332 4593 10367 4627
rect 10401 4593 10436 4627
rect 10470 4593 10505 4627
rect 10539 4593 10574 4627
rect 10608 4593 10643 4627
rect 10677 4593 10712 4627
rect 10746 4593 10781 4627
rect 10815 4593 10850 4627
rect 10884 4593 10919 4627
rect 10953 4593 10987 4627
rect 11021 4593 11055 4627
rect 11089 4593 11123 4627
rect 11157 4593 11191 4627
rect 11225 4593 11259 4627
rect 11293 4593 11327 4627
rect 11361 4593 11395 4627
rect 11429 4593 11463 4627
rect 11497 4593 11531 4627
rect 11565 4593 11599 4627
rect 11633 4593 11667 4627
rect 11701 4593 11735 4627
rect 11769 4593 11803 4627
rect 11837 4593 11871 4627
rect 11905 4593 11939 4627
rect 11973 4593 12007 4627
rect 12041 4593 12075 4627
rect 12109 4593 12143 4627
rect 12177 4593 12211 4627
rect 12245 4593 12279 4627
rect 12313 4593 12347 4627
rect 12381 4593 12415 4627
rect 12449 4593 12483 4627
rect 12517 4593 12551 4627
rect 12585 4593 12619 4627
rect 12653 4593 12687 4627
rect 12721 4593 12755 4627
rect 12789 4593 12823 4627
rect 12857 4593 12891 4627
rect 12925 4593 12959 4627
rect 12993 4593 13027 4627
rect 13061 4593 13095 4627
rect 13129 4593 13163 4627
rect 13197 4593 13231 4627
rect 13265 4593 13367 4627
rect 3442 4588 3510 4593
rect 3340 4587 3510 4588
rect 3374 4557 3510 4587
rect 3374 4553 3476 4557
rect 3340 4549 3476 4553
rect 3340 4517 3408 4549
rect 3374 4515 3408 4517
rect 3442 4523 3476 4549
rect 3442 4515 3510 4523
rect 3374 4487 3510 4515
rect 3374 4483 3476 4487
rect 3340 4476 3476 4483
rect 3340 4447 3408 4476
rect 3374 4442 3408 4447
rect 3442 4453 3476 4476
rect 3442 4442 3510 4453
rect 3374 4417 3510 4442
rect 3374 4413 3476 4417
rect 3340 4403 3476 4413
rect 3340 4377 3408 4403
rect 3374 4369 3408 4377
rect 3442 4383 3476 4403
rect 3442 4369 3510 4383
rect 3374 4347 3510 4369
rect 3374 4343 3476 4347
rect 3340 4330 3476 4343
rect 3340 4307 3408 4330
rect 3374 4296 3408 4307
rect 3442 4313 3476 4330
rect 3442 4296 3510 4313
rect 3374 4277 3510 4296
rect 3374 4273 3476 4277
rect 3340 4256 3476 4273
rect 3340 4237 3408 4256
rect 3374 4222 3408 4237
rect 3442 4243 3476 4256
rect 3442 4222 3510 4243
rect 3374 4207 3510 4222
rect 3374 4203 3476 4207
rect 3340 4182 3476 4203
rect 3340 4167 3408 4182
rect 3374 4148 3408 4167
rect 3442 4173 3476 4182
rect 3442 4148 3510 4173
rect 3374 4136 3510 4148
rect 3374 4133 3476 4136
rect 3340 4108 3476 4133
rect 3340 4096 3408 4108
rect 3374 4074 3408 4096
rect 3442 4102 3476 4108
rect 3442 4074 3510 4102
rect 3374 4065 3510 4074
rect 3374 4062 3476 4065
rect 3340 4034 3476 4062
rect 3340 4025 3408 4034
rect 3374 4000 3408 4025
rect 3442 4031 3476 4034
rect 3442 4000 3510 4031
rect 3374 3994 3510 4000
rect 3374 3991 3476 3994
rect 3340 3960 3476 3991
rect 3340 3954 3408 3960
rect -25 3920 -1 3954
rect 33 3920 68 3954
rect 102 3920 137 3954
rect 171 3920 206 3954
rect 240 3920 275 3954
rect 309 3920 344 3954
rect 378 3920 413 3954
rect 447 3920 482 3954
rect 516 3920 551 3954
rect 585 3920 620 3954
rect -25 3886 620 3920
rect 3374 3926 3408 3954
rect 3442 3926 3510 3960
rect 3374 3923 3510 3926
rect 3374 3889 3476 3923
rect 3374 3886 3510 3889
rect -25 3852 -1 3886
rect 33 3852 68 3886
rect 102 3852 137 3886
rect 171 3852 206 3886
rect 240 3852 275 3886
rect 309 3852 344 3886
rect 378 3852 413 3886
rect 447 3852 482 3886
rect 516 3852 551 3886
rect 585 3852 620 3886
rect 3442 3852 3510 3886
rect -25 3818 2966 3852
rect -25 3784 -1 3818
rect 33 3784 68 3818
rect 102 3784 137 3818
rect 171 3784 206 3818
rect 240 3784 275 3818
rect 309 3784 344 3818
rect 378 3784 413 3818
rect 447 3784 482 3818
rect 516 3784 551 3818
rect 585 3784 620 3818
rect 654 3784 689 3818
rect 723 3784 758 3818
rect 792 3784 827 3818
rect 861 3784 896 3818
rect 930 3784 965 3818
rect 999 3784 1034 3818
rect 1068 3784 1103 3818
rect 1137 3784 1172 3818
rect 1206 3784 1241 3818
rect 1275 3784 1310 3818
rect 1344 3784 1379 3818
rect 1413 3784 1448 3818
rect 1482 3784 1517 3818
rect 1551 3784 1586 3818
rect 1620 3784 1655 3818
rect 1689 3784 1724 3818
rect 1758 3784 1793 3818
rect 1827 3784 1862 3818
rect 1896 3784 1931 3818
rect 1965 3784 2000 3818
rect 2034 3784 2069 3818
rect 2103 3784 2138 3818
rect 2172 3784 2207 3818
rect 2241 3784 2276 3818
rect 2310 3784 2345 3818
rect 2379 3784 2414 3818
rect 2448 3784 2483 3818
rect 2517 3784 2552 3818
rect 2586 3784 2621 3818
rect 2655 3784 2690 3818
rect 2724 3784 2759 3818
rect 2793 3784 2828 3818
rect 2862 3784 2897 3818
rect 2931 3784 2966 3818
rect 3408 3818 3476 3852
rect 3408 3784 3510 3818
rect 19091 2247 19193 2271
rect 19125 2213 19159 2247
rect 19091 2176 19193 2213
rect 19125 2142 19159 2176
rect 19091 2105 19193 2142
rect 19125 2071 19159 2105
rect 19091 2034 19193 2071
rect 19125 2000 19159 2034
rect 19091 1963 19193 2000
rect 19125 1929 19159 1963
rect 19091 1892 19193 1929
rect 19125 1858 19159 1892
rect 19091 1821 19193 1858
rect 19125 1787 19159 1821
rect 19091 1750 19193 1787
rect 19125 1716 19159 1750
rect 19091 1679 19193 1716
rect 19125 1645 19159 1679
rect 19091 1608 19193 1645
rect 19125 1574 19159 1608
rect 19091 1537 19193 1574
rect 19125 1503 19159 1537
rect 19091 1466 19193 1503
rect 19125 1432 19159 1466
rect 19091 1396 19193 1432
rect 19125 1362 19159 1396
rect 19091 1326 19193 1362
rect 19125 1292 19159 1326
rect 19091 1256 19193 1292
rect 19125 1222 19159 1256
rect 19091 1186 19193 1222
rect 19125 1152 19159 1186
rect 19091 1116 19193 1152
rect 19125 1082 19159 1116
rect 19091 1046 19193 1082
rect 19125 1012 19159 1046
rect 19091 976 19193 1012
rect 19125 942 19159 976
rect 19091 918 19193 942
<< mvpsubdiffcont >>
rect 13058 2979 13092 3013
rect 13127 2979 13161 3013
rect 13196 2979 13230 3013
rect 13265 2979 13299 3013
rect 13334 2979 13368 3013
rect 13403 2979 13437 3013
rect 13472 2979 13506 3013
rect 13541 2979 13575 3013
rect 13610 2979 13644 3013
rect 13679 2979 13713 3013
rect 13748 2979 13782 3013
rect 13817 2979 13851 3013
rect 13886 2979 13920 3013
rect 13955 2979 13989 3013
rect 14024 2979 14058 3013
rect 14093 2979 14127 3013
rect 14162 2979 14196 3013
rect 14231 2979 14265 3013
rect 14299 2979 14333 3013
rect 14367 2979 14401 3013
rect 14435 2979 14469 3013
rect 14503 2979 14537 3013
rect 14571 2979 14605 3013
rect 14639 2979 14673 3013
rect 14707 2979 14741 3013
rect 14775 2979 14809 3013
rect 14843 2979 14877 3013
rect 14911 2979 14945 3013
rect 14979 2979 15013 3013
rect 15047 2979 15081 3013
rect 15115 2979 15149 3013
rect 15183 2979 15217 3013
rect 15251 2979 15285 3013
rect 15319 2979 15353 3013
rect 15387 2979 15421 3013
rect 15455 2979 15489 3013
rect 15523 2979 15557 3013
rect 15591 2979 15625 3013
rect 15659 2979 15693 3013
rect 15727 2979 15761 3013
rect 15795 2979 15829 3013
rect 15863 2979 15897 3013
rect 15931 2979 15965 3013
rect 15999 2979 16033 3013
rect 16067 2979 16101 3013
rect 16135 2979 16169 3013
rect 16203 2979 16237 3013
rect 16271 2979 16305 3013
rect 16339 2979 16373 3013
rect 16407 2979 16441 3013
rect 16475 2979 16509 3013
rect 16543 2979 16577 3013
rect 16611 2979 16645 3013
rect 16679 2979 16713 3013
rect 16747 2979 16781 3013
rect 16815 2979 16849 3013
rect 16883 2979 16917 3013
rect 16951 2979 16985 3013
rect 17019 2979 17053 3013
rect 17087 2979 17121 3013
rect 17155 2979 17189 3013
rect 17223 2979 17257 3013
rect 17291 2979 17325 3013
rect 17359 2979 17393 3013
rect 17427 2979 17461 3013
rect 17495 2979 17529 3013
rect 17563 2979 17597 3013
rect 17631 2979 17665 3013
rect 17699 2979 17733 3013
rect 17767 2979 17801 3013
rect 17835 2979 17869 3013
rect 17903 2979 17937 3013
rect 17971 2979 18005 3013
rect 18039 2979 19025 3013
rect 18067 2945 19025 2979
rect 19093 2945 19127 2979
rect 15169 2911 15203 2945
rect 15238 2911 15272 2945
rect 15307 2911 15341 2945
rect 15376 2911 15410 2945
rect 15445 2911 15479 2945
rect 15514 2911 15548 2945
rect 15583 2911 15617 2945
rect 15652 2911 15686 2945
rect 15721 2911 15755 2945
rect 15790 2911 15824 2945
rect 15859 2911 15893 2945
rect 15928 2911 15962 2945
rect 15997 2911 16031 2945
rect 16066 2911 16100 2945
rect 16135 2911 16169 2945
rect 16204 2911 16238 2945
rect 16273 2911 16307 2945
rect 16342 2911 16376 2945
rect 16411 2911 16445 2945
rect 16480 2911 16514 2945
rect 16549 2911 16583 2945
rect 16618 2911 16652 2945
rect 16687 2911 16721 2945
rect 16756 2911 16790 2945
rect 16825 2911 16859 2945
rect 16894 2911 16928 2945
rect 16963 2911 16997 2945
rect 17032 2911 17066 2945
rect 17101 2911 17135 2945
rect 17170 2911 17204 2945
rect 17239 2911 17273 2945
rect 17308 2911 17342 2945
rect 17377 2911 17411 2945
rect 17446 2911 17480 2945
rect 17515 2911 17549 2945
rect 17584 2911 17618 2945
rect 17653 2911 17687 2945
rect 17722 2911 17756 2945
rect 17791 2911 17825 2945
rect 17860 2911 17894 2945
rect 17929 2911 17963 2945
rect 17998 2911 18032 2945
rect 13058 2877 13092 2911
rect 13127 2877 13161 2911
rect 13196 2877 13230 2911
rect 13265 2877 13299 2911
rect 13334 2877 13368 2911
rect 13403 2877 13437 2911
rect 13472 2877 13506 2911
rect 13541 2877 13575 2911
rect 13610 2877 13644 2911
rect 13679 2877 13713 2911
rect 13748 2877 13782 2911
rect 13817 2877 13851 2911
rect 13886 2877 13920 2911
rect 13954 2877 13988 2911
rect 14022 2877 14056 2911
rect 14090 2877 14124 2911
rect 14158 2877 14192 2911
rect 14226 2877 14260 2911
rect 14294 2877 14328 2911
rect 14362 2877 14396 2911
rect 14430 2877 14464 2911
rect 14498 2877 14532 2911
rect 14566 2877 14600 2911
rect 14634 2877 14668 2911
rect 14702 2877 14736 2911
rect 14770 2877 14804 2911
rect 14838 2877 14872 2911
rect 14906 2877 14940 2911
rect 14974 2877 15008 2911
rect 15042 2877 15076 2911
rect 13058 2775 13092 2809
rect 13126 2775 13160 2809
rect 13194 2775 13228 2809
rect 13262 2775 13296 2809
rect 13330 2775 13364 2809
rect 13398 2775 13432 2809
rect 13466 2775 13500 2809
rect 15169 2843 15203 2877
rect 15238 2843 15272 2877
rect 15307 2843 15341 2877
rect 15376 2843 15410 2877
rect 15445 2843 15479 2877
rect 15514 2843 15548 2877
rect 15583 2843 15617 2877
rect 15652 2843 15686 2877
rect 15721 2843 15755 2877
rect 15790 2843 15824 2877
rect 15859 2843 15893 2877
rect 15928 2843 15962 2877
rect 15997 2843 16031 2877
rect 16066 2843 16100 2877
rect 16135 2843 16169 2877
rect 16204 2843 16238 2877
rect 16273 2843 16307 2877
rect 16342 2843 16376 2877
rect 16411 2843 16445 2877
rect 16480 2843 16514 2877
rect 16549 2843 16583 2877
rect 16618 2843 16652 2877
rect 16687 2843 16721 2877
rect 16756 2843 16790 2877
rect 16825 2843 16859 2877
rect 16894 2843 16928 2877
rect 16963 2843 16997 2877
rect 17032 2843 17066 2877
rect 17101 2843 17135 2877
rect 17170 2843 17204 2877
rect 17239 2843 17273 2877
rect 17308 2843 17342 2877
rect 17377 2843 17411 2877
rect 17446 2843 17480 2877
rect 17515 2843 17549 2877
rect 17584 2843 17618 2877
rect 17653 2843 17687 2877
rect 17722 2843 17756 2877
rect 17791 2843 17825 2877
rect 17860 2843 17894 2877
rect 17929 2843 17963 2877
rect 17998 2843 18032 2877
rect 18067 2843 19053 2945
rect 19093 2876 19127 2910
rect 19093 2807 19127 2841
rect 13058 2705 13092 2739
rect 13126 2705 13160 2739
rect 13194 2705 13228 2739
rect 13262 2705 13296 2739
rect 13330 2705 13364 2739
rect 13398 2705 13432 2739
rect 13466 2705 13500 2739
rect 13058 2635 13092 2669
rect 13126 2635 13160 2669
rect 13194 2635 13228 2669
rect 13262 2635 13296 2669
rect 13330 2635 13364 2669
rect 13398 2635 13432 2669
rect 13466 2635 13500 2669
rect 13058 2565 13092 2599
rect 13126 2565 13160 2599
rect 13194 2565 13228 2599
rect 13262 2565 13296 2599
rect 13330 2565 13364 2599
rect 13398 2565 13432 2599
rect 13466 2565 13500 2599
rect 13058 2495 13092 2529
rect 13126 2495 13160 2529
rect 13194 2495 13228 2529
rect 13262 2495 13296 2529
rect 13330 2495 13364 2529
rect 13398 2495 13432 2529
rect 13466 2495 13500 2529
rect 13058 2426 13092 2460
rect 13126 2426 13160 2460
rect 13194 2426 13228 2460
rect 13262 2426 13296 2460
rect 13330 2426 13364 2460
rect 13398 2426 13432 2460
rect 13466 2426 13500 2460
rect 19093 2738 19127 2772
rect 19093 2669 19127 2703
rect 19093 2600 19127 2634
rect 19093 2531 19127 2565
rect 19093 2462 19127 2496
rect 13058 2357 13092 2391
rect 13126 2357 13160 2391
rect 13194 2357 13228 2391
rect 13262 2357 13296 2391
rect 13330 2357 13364 2391
rect 13398 2357 13432 2391
rect 13466 2357 13500 2391
rect 13058 2288 13092 2322
rect 13126 2288 13160 2322
rect 13194 2288 13228 2322
rect 13262 2288 13296 2322
rect 13330 2288 13364 2322
rect 13398 2288 13432 2322
rect 13466 2288 13500 2322
rect 13058 2219 13092 2253
rect 13126 2219 13160 2253
rect 13194 2219 13228 2253
rect 13262 2219 13296 2253
rect 13330 2219 13364 2253
rect 13398 2219 13432 2253
rect 13466 2219 13500 2253
rect 13058 2150 13092 2184
rect 13126 2150 13160 2184
rect 13194 2150 13228 2184
rect 13262 2150 13296 2184
rect 13330 2150 13364 2184
rect 13398 2150 13432 2184
rect 13466 2150 13500 2184
rect 13058 2081 13092 2115
rect 13126 2081 13160 2115
rect 13194 2081 13228 2115
rect 13262 2081 13296 2115
rect 13330 2081 13364 2115
rect 13398 2081 13432 2115
rect 13466 2081 13500 2115
rect 13058 2012 13092 2046
rect 13126 2012 13160 2046
rect 13194 2012 13228 2046
rect 13262 2012 13296 2046
rect 13330 2012 13364 2046
rect 13398 2012 13432 2046
rect 13466 2012 13500 2046
rect 13058 1943 13092 1977
rect 13126 1943 13160 1977
rect 13194 1943 13228 1977
rect 13262 1943 13296 1977
rect 13330 1943 13364 1977
rect 13398 1943 13432 1977
rect 13466 1943 13500 1977
rect 13058 1874 13092 1908
rect 13126 1874 13160 1908
rect 13194 1874 13228 1908
rect 13262 1874 13296 1908
rect 13330 1874 13364 1908
rect 13398 1874 13432 1908
rect 13466 1874 13500 1908
rect 13058 1805 13092 1839
rect 13126 1805 13160 1839
rect 13194 1805 13228 1839
rect 13262 1805 13296 1839
rect 13330 1805 13364 1839
rect 13398 1805 13432 1839
rect 13466 1805 13500 1839
rect 13058 1736 13092 1770
rect 13126 1736 13160 1770
rect 13194 1736 13228 1770
rect 13262 1736 13296 1770
rect 13330 1736 13364 1770
rect 13398 1736 13432 1770
rect 13466 1736 13500 1770
rect 13058 1667 13092 1701
rect 13126 1667 13160 1701
rect 13194 1667 13228 1701
rect 13262 1667 13296 1701
rect 13330 1667 13364 1701
rect 13398 1667 13432 1701
rect 13466 1667 13500 1701
rect 13058 1598 13092 1632
rect 13126 1598 13160 1632
rect 13194 1598 13228 1632
rect 13262 1598 13296 1632
rect 13330 1598 13364 1632
rect 13398 1598 13432 1632
rect 13466 1598 13500 1632
rect 13058 1529 13092 1563
rect 13126 1529 13160 1563
rect 13194 1529 13228 1563
rect 13262 1529 13296 1563
rect 13330 1529 13364 1563
rect 13398 1529 13432 1563
rect 13466 1529 13500 1563
rect 10653 1392 10687 1426
rect 10722 1392 10756 1426
rect 10791 1392 10825 1426
rect 10860 1392 10894 1426
rect 10929 1392 10963 1426
rect 10998 1392 11032 1426
rect 11067 1392 11101 1426
rect 11136 1392 11170 1426
rect 11205 1392 11239 1426
rect 11274 1392 11308 1426
rect 11343 1392 11377 1426
rect 11412 1392 11446 1426
rect 11481 1392 11515 1426
rect 11550 1392 11584 1426
rect 11619 1392 11653 1426
rect 11688 1392 11722 1426
rect 11757 1392 11791 1426
rect 11826 1392 11860 1426
rect 11895 1392 11929 1426
rect 11964 1392 11998 1426
rect 12033 1392 12067 1426
rect 12102 1392 12136 1426
rect 12171 1392 12205 1426
rect 12240 1392 12274 1426
rect 12309 1392 12343 1426
rect 12378 1392 12412 1426
rect 12447 1392 12481 1426
rect 12516 1392 12550 1426
rect 12585 1392 12619 1426
rect 12653 1392 12687 1426
rect 12721 1392 12755 1426
rect 12789 1392 12823 1426
rect 12857 1392 12891 1426
rect 12925 1392 12959 1426
rect 12993 1392 13027 1426
rect 13058 1392 13231 1494
rect 13262 1460 13500 1494
rect 13279 1426 13500 1460
rect 13279 1392 13517 1426
rect 13551 1392 13585 1426
rect 19052 706 19086 740
rect 19052 633 19086 667
rect 19052 560 19086 594
rect 19052 488 19086 522
rect 10619 394 10653 428
rect 10619 304 10653 338
rect 19052 416 19086 450
rect 19052 344 19086 378
rect 10721 294 10755 328
rect 10790 294 10824 328
rect 10859 294 10893 328
rect 10928 294 10962 328
rect 10997 294 11031 328
rect 11066 294 11100 328
rect 11135 294 11169 328
rect 11204 294 11238 328
rect 11273 294 11307 328
rect 11342 294 11376 328
rect 11411 294 11445 328
rect 11480 294 11514 328
rect 11549 294 11583 328
rect 11618 294 11652 328
rect 11687 294 11721 328
rect 11756 294 11790 328
rect 11825 294 11859 328
rect 11894 294 11928 328
rect 11963 294 11997 328
rect 12032 294 12066 328
rect 12101 294 12135 328
rect 12170 294 12204 328
rect 12239 294 12273 328
rect 12308 294 12342 328
rect 12377 294 12411 328
rect 12446 294 12480 328
rect 12515 294 12549 328
rect 12584 294 12618 328
rect 12653 294 12687 328
rect 12722 294 12756 328
rect 12791 294 12825 328
rect 12860 294 12894 328
rect 12929 294 12963 328
rect 12998 294 13032 328
rect 10619 214 10653 248
rect 10721 226 10755 260
rect 10790 226 10824 260
rect 10859 226 10893 260
rect 10928 226 10962 260
rect 10997 226 11031 260
rect 11066 226 11100 260
rect 11135 226 11169 260
rect 11204 226 11238 260
rect 11273 226 11307 260
rect 11342 226 11376 260
rect 11411 226 11445 260
rect 11480 226 11514 260
rect 11549 226 11583 260
rect 11618 226 11652 260
rect 11687 226 11721 260
rect 11756 226 11790 260
rect 11825 226 11859 260
rect 11894 226 11928 260
rect 11963 226 11997 260
rect 12032 226 12066 260
rect 12101 226 12135 260
rect 12170 226 12204 260
rect 12239 226 12273 260
rect 12308 226 12342 260
rect 12377 226 12411 260
rect 12446 226 12480 260
rect 12515 226 12549 260
rect 12584 226 12618 260
rect 12653 226 12687 260
rect 12722 226 12756 260
rect 12791 226 12825 260
rect 12860 226 12894 260
rect 12929 226 12963 260
rect 12998 226 13032 260
rect 10721 158 10755 192
rect 10790 158 10824 192
rect 10859 158 10893 192
rect 10928 158 10962 192
rect 10997 158 11031 192
rect 11066 158 11100 192
rect 11135 158 11169 192
rect 11204 158 11238 192
rect 11273 158 11307 192
rect 11342 158 11376 192
rect 11411 158 11445 192
rect 11480 158 11514 192
rect 11549 158 11583 192
rect 11618 158 11652 192
rect 11687 158 11721 192
rect 11756 158 11790 192
rect 11825 158 11859 192
rect 11894 158 11928 192
rect 11963 158 11997 192
rect 12032 158 12066 192
rect 12101 158 12135 192
rect 12170 158 12204 192
rect 12239 158 12273 192
rect 12308 158 12342 192
rect 12377 158 12411 192
rect 12446 158 12480 192
rect 12515 158 12549 192
rect 12584 158 12618 192
rect 12653 158 12687 192
rect 12722 158 12756 192
rect 12791 158 12825 192
rect 12860 158 12894 192
rect 12929 158 12963 192
rect 12998 158 13032 192
rect 10619 124 10653 158
rect 13067 124 15073 328
rect 15171 260 15205 294
rect 15240 260 15274 294
rect 15309 260 15343 294
rect 15378 260 15412 294
rect 15447 260 15481 294
rect 15516 260 15550 294
rect 15585 260 15619 294
rect 15654 260 15688 294
rect 15723 260 15757 294
rect 15792 260 15826 294
rect 15861 260 15895 294
rect 15930 260 15964 294
rect 15999 260 16033 294
rect 16068 260 16102 294
rect 16137 260 16171 294
rect 16206 260 16240 294
rect 16275 260 16309 294
rect 16344 260 16378 294
rect 16413 260 16447 294
rect 16482 260 16516 294
rect 16551 260 16585 294
rect 16620 260 16654 294
rect 16689 260 16723 294
rect 16758 260 16792 294
rect 16827 260 16861 294
rect 16896 260 16930 294
rect 16965 260 16999 294
rect 17034 260 17068 294
rect 17103 260 17137 294
rect 17172 260 17206 294
rect 17241 260 17275 294
rect 17310 260 17344 294
rect 17379 260 17413 294
rect 17448 260 17482 294
rect 17517 260 17551 294
rect 17586 260 17620 294
rect 17655 260 17689 294
rect 17724 260 17758 294
rect 17793 260 17827 294
rect 17862 260 17896 294
rect 17931 260 17965 294
rect 18000 260 18034 294
rect 18069 260 18103 294
rect 18138 260 18172 294
rect 18208 260 18242 294
rect 18278 260 18312 294
rect 18348 260 18382 294
rect 18418 260 18452 294
rect 18488 260 18522 294
rect 18558 260 18592 294
rect 18628 260 18662 294
rect 18698 260 18732 294
rect 18768 260 18802 294
rect 18838 260 18872 294
rect 18908 260 18942 294
rect 18978 260 19012 294
rect 19052 272 19086 306
rect 15171 192 15205 226
rect 15240 192 15274 226
rect 15309 192 15343 226
rect 15378 192 15412 226
rect 15447 192 15481 226
rect 15516 192 15550 226
rect 15585 192 15619 226
rect 15654 192 15688 226
rect 15723 192 15757 226
rect 15792 192 15826 226
rect 15861 192 15895 226
rect 15930 192 15964 226
rect 15999 192 16033 226
rect 16068 192 16102 226
rect 16137 192 16171 226
rect 16206 192 16240 226
rect 16275 192 16309 226
rect 16344 192 16378 226
rect 16413 192 16447 226
rect 16482 192 16516 226
rect 16551 192 16585 226
rect 16620 192 16654 226
rect 16689 192 16723 226
rect 16758 192 16792 226
rect 16827 192 16861 226
rect 16896 192 16930 226
rect 16965 192 16999 226
rect 17034 192 17068 226
rect 17103 192 17137 226
rect 17172 192 17206 226
rect 17241 192 17275 226
rect 17310 192 17344 226
rect 17379 192 17413 226
rect 17448 192 17482 226
rect 17517 192 17551 226
rect 17586 192 17620 226
rect 17655 192 17689 226
rect 17724 192 17758 226
rect 17793 192 17827 226
rect 17862 192 17896 226
rect 17931 192 17965 226
rect 18000 192 18034 226
rect 18069 192 18103 226
rect 18138 192 18172 226
rect 18208 192 18242 226
rect 18278 192 18312 226
rect 18348 192 18382 226
rect 18418 192 18452 226
rect 18488 192 18522 226
rect 18558 192 18592 226
rect 18628 192 18662 226
rect 18698 192 18732 226
rect 18768 192 18802 226
rect 18838 192 18872 226
rect 18908 192 18942 226
rect 18978 192 19012 226
rect 19052 200 19086 234
rect 10721 90 10755 124
rect 10789 90 10823 124
rect 10857 90 10891 124
rect 10925 90 10959 124
rect 10993 90 11027 124
rect 11061 90 11095 124
rect 11129 90 11163 124
rect 11197 90 11231 124
rect 11265 90 11299 124
rect 11333 90 11367 124
rect 11401 90 11435 124
rect 11469 90 11503 124
rect 11537 90 11571 124
rect 11605 90 11639 124
rect 11673 90 11707 124
rect 11741 90 11775 124
rect 11809 90 11843 124
rect 11877 90 11911 124
rect 11945 90 11979 124
rect 12013 90 12047 124
rect 12081 90 12115 124
rect 12149 90 12183 124
rect 12217 90 12251 124
rect 12285 90 12319 124
rect 12353 90 12387 124
rect 12421 90 12455 124
rect 12489 90 12523 124
rect 12557 90 12591 124
rect 12625 90 12659 124
rect 12693 90 12727 124
rect 12761 90 12795 124
rect 12829 90 12863 124
rect 12897 90 12931 124
rect 12965 90 12999 124
rect 13033 90 15107 124
rect 15141 90 15175 124
rect 15209 90 15243 124
rect 15277 90 15311 124
rect 15345 90 15379 124
rect 15413 90 15447 124
rect 15481 90 15515 124
rect 15549 90 15583 124
rect 15617 90 15651 124
rect 15685 90 15719 124
rect 15753 90 15787 124
rect 15821 90 15855 124
rect 15889 90 15923 124
rect 15957 90 15991 124
rect 16025 90 16059 124
rect 16093 90 16127 124
rect 16161 90 16195 124
rect 16229 90 16263 124
rect 16297 90 16331 124
rect 16365 90 16399 124
rect 16433 90 16467 124
rect 16501 90 16535 124
rect 16569 90 16603 124
rect 16637 90 16671 124
rect 16705 90 16739 124
rect 16773 90 16807 124
rect 16841 90 16875 124
rect 16909 90 16943 124
rect 16977 90 17011 124
rect 17045 90 17079 124
rect 17113 90 17147 124
rect 17181 90 17215 124
rect 17249 90 17283 124
rect 17317 90 17351 124
rect 17385 90 17419 124
rect 17453 90 17487 124
rect 17521 90 17555 124
rect 17589 90 17623 124
rect 17657 90 17691 124
rect 17725 90 17759 124
rect 17793 90 17827 124
rect 17861 90 17895 124
rect 17929 90 17963 124
rect 17997 90 18031 124
rect 18065 90 18099 124
rect 18133 90 18167 124
rect 18201 90 18235 124
rect 18269 90 18303 124
rect 18337 90 18371 124
rect 18405 90 18439 124
rect 18473 90 18507 124
rect 18541 90 18575 124
rect 18609 90 18643 124
rect 18677 90 18711 124
rect 18745 90 18779 124
rect 18813 90 18847 124
rect 18881 90 18915 124
rect 18949 90 18983 124
rect 19018 90 19052 124
<< mvnsubdiffcont >>
rect -1 6906 33 6940
rect 68 6906 102 6940
rect 137 6906 171 6940
rect 206 6906 240 6940
rect 275 6906 309 6940
rect 344 6906 378 6940
rect 413 6906 447 6940
rect 482 6906 516 6940
rect 551 6906 585 6940
rect 620 6906 654 6940
rect 689 6906 723 6940
rect 758 6906 792 6940
rect 827 6906 861 6940
rect 896 6906 930 6940
rect 965 6906 999 6940
rect 1034 6906 1068 6940
rect 1103 6906 1137 6940
rect 1172 6906 1206 6940
rect 1241 6906 1275 6940
rect 1310 6906 1344 6940
rect 1379 6906 1413 6940
rect 1448 6906 1482 6940
rect 1517 6906 1551 6940
rect 1586 6906 1620 6940
rect 1655 6906 1689 6940
rect 1724 6906 1758 6940
rect 1793 6906 1827 6940
rect -1 6838 33 6872
rect 68 6838 102 6872
rect 137 6838 171 6872
rect 206 6838 240 6872
rect 275 6838 309 6872
rect 344 6838 378 6872
rect 413 6838 447 6872
rect 482 6838 516 6872
rect 551 6838 585 6872
rect 620 6838 654 6872
rect 689 6838 723 6872
rect 758 6838 792 6872
rect 827 6838 861 6872
rect 896 6838 930 6872
rect 965 6838 999 6872
rect 1034 6838 1068 6872
rect 1103 6838 1137 6872
rect 1172 6838 1206 6872
rect 1241 6838 1275 6872
rect 1310 6838 1344 6872
rect 1379 6838 1413 6872
rect 1448 6838 1482 6872
rect 1517 6838 1551 6872
rect 1586 6838 1620 6872
rect 1655 6838 1689 6872
rect 1724 6838 1758 6872
rect 1793 6838 1827 6872
rect -1 6770 33 6804
rect 68 6770 102 6804
rect 137 6770 171 6804
rect 206 6770 240 6804
rect 275 6770 309 6804
rect 344 6770 378 6804
rect 413 6770 447 6804
rect 482 6770 516 6804
rect 551 6770 585 6804
rect 620 6770 654 6804
rect 689 6770 723 6804
rect 758 6770 792 6804
rect 827 6770 861 6804
rect 896 6770 930 6804
rect 965 6770 999 6804
rect 1034 6770 1068 6804
rect 1103 6770 1137 6804
rect 1172 6770 1206 6804
rect 1241 6770 1275 6804
rect 1310 6770 1344 6804
rect 1379 6770 1413 6804
rect 1448 6770 1482 6804
rect 1517 6770 1551 6804
rect 1586 6770 1620 6804
rect 1655 6770 1689 6804
rect 1724 6770 1758 6804
rect 1793 6770 1827 6804
rect 1862 6770 10056 6940
rect 10090 6906 10124 6940
rect 10158 6906 10192 6940
rect 10226 6906 10260 6940
rect 10294 6906 10328 6940
rect 10362 6906 10396 6940
rect 10430 6906 10464 6940
rect 10498 6906 10532 6940
rect 10566 6906 10600 6940
rect 10634 6906 10668 6940
rect 10702 6906 10736 6940
rect 10770 6906 10804 6940
rect 10838 6906 10872 6940
rect 10906 6906 10940 6940
rect 10974 6906 11008 6940
rect 11042 6906 11076 6940
rect 11110 6906 11144 6940
rect 11178 6906 11212 6940
rect 11246 6906 11280 6940
rect 11314 6906 11348 6940
rect 11382 6906 11416 6940
rect 11450 6906 11484 6940
rect 11518 6906 11552 6940
rect 11586 6906 11620 6940
rect 11654 6906 11688 6940
rect 11722 6906 11756 6940
rect 11790 6906 11824 6940
rect 11858 6906 11892 6940
rect 11926 6906 11960 6940
rect 11994 6906 12028 6940
rect 12062 6906 12096 6940
rect 12130 6906 12164 6940
rect 12198 6906 12232 6940
rect 12266 6906 12300 6940
rect 12334 6906 12368 6940
rect 12402 6906 12436 6940
rect 12471 6906 12505 6940
rect 12540 6906 12574 6940
rect 12609 6906 12643 6940
rect 12678 6906 12712 6940
rect 12747 6906 12781 6940
rect 12816 6906 12850 6940
rect 12885 6906 12919 6940
rect 12954 6906 12988 6940
rect 13023 6906 13057 6940
rect 13092 6906 13126 6940
rect 13161 6906 13195 6940
rect 13230 6906 13264 6940
rect 13299 6906 13333 6940
rect 10091 6838 10125 6872
rect 10160 6838 10194 6872
rect 10229 6838 10263 6872
rect 10298 6838 10332 6872
rect 10367 6838 10401 6872
rect 10436 6838 10470 6872
rect 10505 6838 10539 6872
rect 10574 6838 10608 6872
rect 10643 6838 10677 6872
rect 10712 6838 10746 6872
rect 10781 6838 10815 6872
rect 10850 6838 10884 6872
rect 10919 6838 10953 6872
rect 10988 6838 11022 6872
rect 11057 6838 11091 6872
rect 11126 6838 11160 6872
rect 11195 6838 11229 6872
rect 11264 6838 11298 6872
rect 11333 6838 11367 6872
rect 11402 6838 11436 6872
rect 11471 6838 11505 6872
rect 11540 6838 11574 6872
rect 11609 6838 11643 6872
rect 11678 6838 11712 6872
rect 11747 6838 11781 6872
rect 11816 6838 11850 6872
rect 11885 6838 11919 6872
rect 11954 6838 11988 6872
rect 12023 6838 12057 6872
rect 12092 6838 12126 6872
rect 12161 6838 12195 6872
rect 12230 6838 12264 6872
rect 12299 6838 12333 6872
rect 12368 6838 12402 6872
rect 12437 6838 12471 6872
rect 12506 6838 12540 6872
rect 12575 6838 12609 6872
rect 12644 6838 12678 6872
rect 12713 6838 12747 6872
rect 12782 6838 12816 6872
rect 12851 6838 12885 6872
rect 12920 6838 12954 6872
rect 12989 6838 13023 6872
rect 13058 6838 13092 6872
rect 13127 6838 13161 6872
rect 13196 6838 13230 6872
rect 13265 6838 13299 6872
rect 13265 6804 13367 6838
rect 10091 6770 10125 6804
rect 10160 6770 10194 6804
rect 10229 6770 10263 6804
rect 10298 6770 10332 6804
rect 10367 6770 10401 6804
rect 10436 6770 10470 6804
rect 10505 6770 10539 6804
rect 10574 6770 10608 6804
rect 10643 6770 10677 6804
rect 10712 6770 10746 6804
rect 10781 6770 10815 6804
rect 10850 6770 10884 6804
rect 10919 6770 10953 6804
rect 10988 6770 11022 6804
rect 11057 6770 11091 6804
rect 11126 6770 11160 6804
rect 11195 6770 11229 6804
rect 11264 6770 11298 6804
rect 11333 6770 11367 6804
rect 11402 6770 11436 6804
rect 11471 6770 11505 6804
rect 11540 6770 11574 6804
rect 11609 6770 11643 6804
rect 11678 6770 11712 6804
rect 11747 6770 11781 6804
rect 11816 6770 11850 6804
rect 11885 6770 11919 6804
rect 11954 6770 11988 6804
rect 12023 6770 12057 6804
rect 12092 6770 12126 6804
rect 12161 6770 12195 6804
rect 12230 6770 12264 6804
rect 12299 6770 12333 6804
rect 12368 6770 12402 6804
rect 12437 6770 12471 6804
rect 12506 6770 12540 6804
rect 12575 6770 12609 6804
rect 12644 6770 12678 6804
rect 12713 6770 12747 6804
rect 12782 6770 12816 6804
rect 12851 6770 12885 6804
rect 12920 6770 12954 6804
rect 12989 6770 13023 6804
rect 13058 6770 13092 6804
rect 13127 6770 13161 6804
rect 3373 6694 3407 6728
rect 3441 6694 3475 6728
rect 3509 6694 3543 6728
rect 3577 6694 3611 6728
rect 3645 6694 3679 6728
rect 3713 6694 3747 6728
rect 3781 6694 3815 6728
rect 3849 6694 3883 6728
rect 3917 6694 3951 6728
rect 3985 6694 4019 6728
rect 4053 6694 4087 6728
rect 4121 6694 4155 6728
rect 4189 6694 4223 6728
rect 4257 6694 4291 6728
rect 4325 6694 4359 6728
rect 4393 6694 4427 6728
rect 4461 6694 4495 6728
rect 4529 6694 4563 6728
rect 4597 6694 4631 6728
rect 4665 6694 4699 6728
rect 4733 6694 4767 6728
rect 4801 6694 4835 6728
rect 4869 6694 4903 6728
rect 4937 6694 4971 6728
rect 5005 6694 5039 6728
rect 5073 6694 5107 6728
rect 5180 6661 5214 6695
rect 5248 6661 5282 6695
rect 5316 6661 5350 6695
rect 5384 6661 5418 6695
rect 5452 6661 5486 6695
rect 5520 6661 5554 6695
rect 3373 6624 3407 6658
rect 3441 6624 3475 6658
rect 3509 6624 3543 6658
rect 3577 6624 3611 6658
rect 3645 6624 3679 6658
rect 3713 6624 3747 6658
rect 3781 6624 3815 6658
rect 3849 6624 3883 6658
rect 3917 6624 3951 6658
rect 3985 6624 4019 6658
rect 4053 6624 4087 6658
rect 4121 6624 4155 6658
rect 4189 6624 4223 6658
rect 4257 6624 4291 6658
rect 4325 6624 4359 6658
rect 4393 6624 4427 6658
rect 4461 6624 4495 6658
rect 4529 6624 4563 6658
rect 4597 6624 4631 6658
rect 4665 6624 4699 6658
rect 4733 6624 4767 6658
rect 4801 6624 4835 6658
rect 4869 6624 4903 6658
rect 4937 6624 4971 6658
rect 5005 6624 5039 6658
rect 5073 6624 5107 6658
rect 5180 6591 5214 6625
rect 5248 6591 5282 6625
rect 5316 6591 5350 6625
rect 5384 6591 5418 6625
rect 5452 6591 5486 6625
rect 5520 6591 5554 6625
rect 6781 6702 6815 6736
rect 6781 6629 6815 6663
rect 3373 6554 3407 6588
rect 3441 6554 3475 6588
rect 3509 6554 3543 6588
rect 3577 6554 3611 6588
rect 3645 6554 3679 6588
rect 3713 6554 3747 6588
rect 3781 6554 3815 6588
rect 3849 6554 3883 6588
rect 3917 6554 3951 6588
rect 3985 6554 4019 6588
rect 4053 6554 4087 6588
rect 4121 6554 4155 6588
rect 4189 6554 4223 6588
rect 4257 6554 4291 6588
rect 4325 6554 4359 6588
rect 4393 6554 4427 6588
rect 4461 6554 4495 6588
rect 4529 6554 4563 6588
rect 4597 6554 4631 6588
rect 4665 6554 4699 6588
rect 4733 6554 4767 6588
rect 4801 6554 4835 6588
rect 4869 6554 4903 6588
rect 4937 6554 4971 6588
rect 5005 6554 5039 6588
rect 5073 6554 5107 6588
rect 5180 6522 5214 6556
rect 5248 6522 5282 6556
rect 5316 6522 5350 6556
rect 5384 6522 5418 6556
rect 5452 6522 5486 6556
rect 5520 6522 5554 6556
rect 3373 6484 3407 6518
rect 3441 6484 3475 6518
rect 3509 6484 3543 6518
rect 3577 6484 3611 6518
rect 3645 6484 3679 6518
rect 3713 6484 3747 6518
rect 3781 6484 3815 6518
rect 3849 6484 3883 6518
rect 3917 6484 3951 6518
rect 3985 6484 4019 6518
rect 4053 6484 4087 6518
rect 4121 6484 4155 6518
rect 4189 6484 4223 6518
rect 4257 6484 4291 6518
rect 4325 6484 4359 6518
rect 4393 6484 4427 6518
rect 4461 6484 4495 6518
rect 4529 6484 4563 6518
rect 4597 6484 4631 6518
rect 4665 6484 4699 6518
rect 4733 6484 4767 6518
rect 4801 6484 4835 6518
rect 4869 6484 4903 6518
rect 4937 6484 4971 6518
rect 5005 6484 5039 6518
rect 5073 6484 5107 6518
rect 5180 6453 5214 6487
rect 5248 6453 5282 6487
rect 5316 6453 5350 6487
rect 5384 6453 5418 6487
rect 5452 6453 5486 6487
rect 5520 6453 5554 6487
rect 3373 6414 3407 6448
rect 3441 6414 3475 6448
rect 3509 6414 3543 6448
rect 3577 6414 3611 6448
rect 3645 6414 3679 6448
rect 3713 6414 3747 6448
rect 3781 6414 3815 6448
rect 3849 6414 3883 6448
rect 3917 6414 3951 6448
rect 3985 6414 4019 6448
rect 4053 6414 4087 6448
rect 4121 6414 4155 6448
rect 4189 6414 4223 6448
rect 4257 6414 4291 6448
rect 4325 6414 4359 6448
rect 4393 6414 4427 6448
rect 4461 6414 4495 6448
rect 4529 6414 4563 6448
rect 4597 6414 4631 6448
rect 4665 6414 4699 6448
rect 4733 6414 4767 6448
rect 4801 6414 4835 6448
rect 4869 6414 4903 6448
rect 4937 6414 4971 6448
rect 5005 6414 5039 6448
rect 5073 6414 5107 6448
rect 6781 6557 6815 6591
rect 6781 6485 6815 6519
rect 9317 6482 13159 6720
rect 5180 6384 5214 6418
rect 5248 6384 5282 6418
rect 5316 6384 5350 6418
rect 5384 6384 5418 6418
rect 5452 6384 5486 6418
rect 5520 6384 5554 6418
rect 6825 6414 6859 6448
rect 6893 6414 6927 6448
rect 6961 6414 6995 6448
rect 7029 6414 7063 6448
rect 7097 6414 7131 6448
rect 7165 6414 7199 6448
rect 7233 6414 7267 6448
rect 7301 6414 7335 6448
rect 7369 6414 7403 6448
rect 7437 6414 7471 6448
rect 7505 6414 7539 6448
rect 7573 6414 7607 6448
rect 7641 6414 7675 6448
rect 7709 6414 7743 6448
rect 7777 6414 7811 6448
rect 7845 6414 7879 6448
rect 7913 6414 7947 6448
rect 7981 6414 8015 6448
rect 8049 6414 8083 6448
rect 8117 6414 8151 6448
rect 8185 6414 8219 6448
rect 8253 6414 8287 6448
rect 8321 6414 8355 6448
rect 8389 6414 8423 6448
rect 8457 6414 8491 6448
rect 8525 6414 8559 6448
rect 8593 6414 8627 6448
rect 8661 6414 8695 6448
rect 8729 6414 8763 6448
rect 8797 6414 8831 6448
rect 8865 6414 8899 6448
rect 8933 6414 8967 6448
rect 9001 6414 9035 6448
rect 9069 6414 9103 6448
rect 9137 6414 9171 6448
rect 9205 6414 9239 6448
rect 9273 6414 9307 6448
rect 9317 6414 9851 6482
rect 9886 6414 9920 6448
rect 9955 6414 9989 6448
rect 10024 6414 10058 6448
rect 10093 6414 10127 6448
rect 10162 6414 10196 6448
rect 10231 6414 10265 6448
rect 10300 6414 10334 6448
rect 10369 6414 10403 6448
rect 10438 6414 10472 6448
rect 10507 6414 10541 6448
rect 10576 6414 10610 6448
rect 10645 6414 10679 6448
rect 10714 6414 10748 6448
rect 10783 6414 10817 6448
rect 10852 6414 10886 6448
rect 10921 6414 10955 6448
rect 10990 6414 11024 6448
rect 11059 6414 11093 6448
rect 11128 6414 11162 6448
rect 11197 6414 11231 6448
rect 11266 6414 11300 6448
rect 11335 6414 11369 6448
rect 11404 6414 11438 6448
rect 11473 6414 11507 6448
rect 11542 6414 11576 6448
rect 11611 6414 11645 6448
rect 11680 6414 11714 6448
rect 11749 6414 11783 6448
rect 11818 6414 11852 6448
rect 11887 6414 11921 6448
rect 11956 6414 11990 6448
rect 12025 6414 12059 6448
rect 12094 6414 12128 6448
rect 12163 6414 12197 6448
rect 12232 6414 12266 6448
rect 12301 6414 12335 6448
rect 12370 6414 12404 6448
rect 12439 6414 12473 6448
rect 12508 6414 12542 6448
rect 12577 6414 12611 6448
rect 12646 6414 12680 6448
rect 12715 6414 12749 6448
rect 12784 6414 12818 6448
rect 12853 6414 12887 6448
rect 12922 6414 12956 6448
rect 12991 6414 13025 6448
rect 13060 6414 13094 6448
rect 13129 6414 13163 6448
rect 3373 6344 3407 6378
rect 3441 6344 3475 6378
rect 3509 6344 3543 6378
rect 3577 6344 3611 6378
rect 3645 6344 3679 6378
rect 3713 6344 3747 6378
rect 3781 6344 3815 6378
rect 3849 6344 3883 6378
rect 3917 6344 3951 6378
rect 3985 6344 4019 6378
rect 4053 6344 4087 6378
rect 4121 6344 4155 6378
rect 4189 6344 4223 6378
rect 4257 6344 4291 6378
rect 4325 6344 4359 6378
rect 4393 6344 4427 6378
rect 4461 6344 4495 6378
rect 4529 6344 4563 6378
rect 4597 6344 4631 6378
rect 4665 6344 4699 6378
rect 4733 6344 4767 6378
rect 4801 6344 4835 6378
rect 4869 6344 4903 6378
rect 4937 6344 4971 6378
rect 5005 6344 5039 6378
rect 5073 6344 5107 6378
rect 5180 6315 5214 6349
rect 5248 6315 5282 6349
rect 5316 6315 5350 6349
rect 5384 6315 5418 6349
rect 5452 6315 5486 6349
rect 5520 6315 5554 6349
rect 3373 6274 3407 6308
rect 3441 6274 3475 6308
rect 3509 6274 3543 6308
rect 3577 6274 3611 6308
rect 3645 6274 3679 6308
rect 3713 6274 3747 6308
rect 3781 6274 3815 6308
rect 3849 6274 3883 6308
rect 3917 6274 3951 6308
rect 3985 6274 4019 6308
rect 4053 6274 4087 6308
rect 4121 6274 4155 6308
rect 4189 6274 4223 6308
rect 4257 6274 4291 6308
rect 4325 6274 4359 6308
rect 4393 6274 4427 6308
rect 4461 6274 4495 6308
rect 4529 6274 4563 6308
rect 4597 6274 4631 6308
rect 4665 6274 4699 6308
rect 4733 6274 4767 6308
rect 4801 6274 4835 6308
rect 4869 6274 4903 6308
rect 4937 6274 4971 6308
rect 5005 6274 5039 6308
rect 5073 6274 5107 6308
rect 3373 6204 3407 6238
rect 3441 6204 3475 6238
rect 3509 6204 3543 6238
rect 3577 6204 3611 6238
rect 3645 6204 3679 6238
rect 3713 6204 3747 6238
rect 3781 6204 3815 6238
rect 3849 6204 3883 6238
rect 3917 6204 3951 6238
rect 3985 6204 4019 6238
rect 4053 6204 4087 6238
rect 4121 6204 4155 6238
rect 4189 6204 4223 6238
rect 4257 6204 4291 6238
rect 4325 6204 4359 6238
rect 4393 6204 4427 6238
rect 4461 6204 4495 6238
rect 4529 6204 4563 6238
rect 4597 6204 4631 6238
rect 4665 6204 4699 6238
rect 4733 6204 4767 6238
rect 4801 6204 4835 6238
rect 4869 6204 4903 6238
rect 4937 6204 4971 6238
rect 5005 6204 5039 6238
rect 5073 6204 5107 6238
rect 5155 6184 5189 6218
rect 5223 6184 5257 6218
rect 5291 6184 5325 6218
rect 5359 6184 5393 6218
rect 5427 6184 5461 6218
rect 5495 6184 5529 6218
rect 5563 6184 5597 6218
rect 5631 6184 5665 6218
rect 5699 6184 5733 6218
rect 5767 6184 5801 6218
rect 5835 6184 5869 6218
rect 5903 6184 5937 6218
rect 5971 6184 6005 6218
rect 6040 6184 6074 6218
rect 6108 6184 6142 6218
rect 6176 6184 6210 6218
rect 6244 6184 6278 6218
rect 6312 6184 6346 6218
rect 6380 6184 6414 6218
rect 6448 6184 6482 6218
rect 6516 6184 6550 6218
rect 6584 6184 6618 6218
rect 6652 6184 6686 6218
rect 6720 6184 6754 6218
rect 3373 6134 3407 6168
rect 3441 6134 3475 6168
rect 3509 6134 3543 6168
rect 3577 6134 3611 6168
rect 3645 6134 3679 6168
rect 3713 6134 3747 6168
rect 3781 6134 3815 6168
rect 3849 6134 3883 6168
rect 3917 6134 3951 6168
rect 3985 6134 4019 6168
rect 4053 6134 4087 6168
rect 4121 6134 4155 6168
rect 4189 6134 4223 6168
rect 4257 6134 4291 6168
rect 4325 6134 4359 6168
rect 4393 6134 4427 6168
rect 4461 6134 4495 6168
rect 4529 6134 4563 6168
rect 4597 6134 4631 6168
rect 4665 6134 4699 6168
rect 4733 6134 4767 6168
rect 4801 6134 4835 6168
rect 4869 6134 4903 6168
rect 4937 6134 4971 6168
rect 5005 6134 5039 6168
rect 5073 6134 5107 6168
rect 5155 6114 5189 6148
rect 5223 6114 5257 6148
rect 5291 6114 5325 6148
rect 5359 6114 5393 6148
rect 5427 6114 5461 6148
rect 5495 6114 5529 6148
rect 5563 6114 5597 6148
rect 5631 6114 5665 6148
rect 5699 6114 5733 6148
rect 5767 6114 5801 6148
rect 5835 6114 5869 6148
rect 5903 6114 5937 6148
rect 5971 6114 6005 6148
rect 6040 6115 6074 6149
rect 6108 6115 6142 6149
rect 6176 6115 6210 6149
rect 6244 6115 6278 6149
rect 6312 6115 6346 6149
rect 6380 6115 6414 6149
rect 6448 6115 6482 6149
rect 6516 6115 6550 6149
rect 6584 6115 6618 6149
rect 6652 6115 6686 6149
rect 6720 6115 6754 6149
rect 3373 6064 3407 6098
rect 3441 6064 3475 6098
rect 3509 6064 3543 6098
rect 3577 6064 3611 6098
rect 3645 6064 3679 6098
rect 3713 6064 3747 6098
rect 3781 6064 3815 6098
rect 3849 6064 3883 6098
rect 3917 6064 3951 6098
rect 3985 6064 4019 6098
rect 4053 6064 4087 6098
rect 4121 6064 4155 6098
rect 4189 6064 4223 6098
rect 4257 6064 4291 6098
rect 4325 6064 4359 6098
rect 4393 6064 4427 6098
rect 4461 6064 4495 6098
rect 4529 6064 4563 6098
rect 4597 6064 4631 6098
rect 4665 6064 4699 6098
rect 4733 6064 4767 6098
rect 4801 6064 4835 6098
rect 4869 6064 4903 6098
rect 4937 6064 4971 6098
rect 5005 6064 5039 6098
rect 5073 6064 5107 6098
rect 5155 6044 5189 6078
rect 5223 6044 5257 6078
rect 5291 6044 5325 6078
rect 5359 6044 5393 6078
rect 5427 6044 5461 6078
rect 5495 6044 5529 6078
rect 5563 6044 5597 6078
rect 5631 6044 5665 6078
rect 5699 6044 5733 6078
rect 5767 6044 5801 6078
rect 5835 6044 5869 6078
rect 5903 6044 5937 6078
rect 5971 6044 6005 6078
rect 6040 6046 6074 6080
rect 6108 6046 6142 6080
rect 6176 6046 6210 6080
rect 6244 6046 6278 6080
rect 6312 6046 6346 6080
rect 6380 6046 6414 6080
rect 6448 6046 6482 6080
rect 6516 6046 6550 6080
rect 6584 6046 6618 6080
rect 6652 6046 6686 6080
rect 6720 6046 6754 6080
rect 6825 6037 6859 6071
rect 6893 6037 6927 6071
rect 6961 6037 6995 6071
rect 7029 6037 7063 6071
rect 7097 6037 7131 6071
rect 7165 6037 7199 6071
rect 7233 6037 7267 6071
rect 7301 6037 7335 6071
rect 7369 6037 7403 6071
rect 7437 6037 7471 6071
rect 7505 6037 7539 6071
rect 7573 6037 7607 6071
rect 7641 6037 7675 6071
rect 7709 6037 7743 6071
rect 7777 6037 7811 6071
rect 7845 6037 7879 6071
rect 7913 6037 7947 6071
rect 7981 6037 8015 6071
rect 8049 6037 8083 6071
rect 8117 6037 8151 6071
rect 8185 6037 8219 6071
rect 8253 6037 8287 6071
rect 8321 6037 8355 6071
rect 8389 6037 8423 6071
rect 8457 6037 8491 6071
rect 8525 6037 8559 6071
rect 8593 6037 8627 6071
rect 8661 6037 8695 6071
rect 8729 6037 8763 6071
rect 8797 6037 8831 6071
rect 8865 6037 8899 6071
rect 8933 6037 8967 6071
rect 9001 6037 9035 6071
rect 9069 6037 9103 6071
rect 9137 6037 9171 6071
rect 9205 6037 9239 6071
rect 9273 6037 9307 6071
rect 9341 6037 9375 6071
rect 9409 6037 9443 6071
rect 9477 6037 9511 6071
rect 9545 6037 9579 6071
rect 9613 6037 9647 6071
rect 9681 6037 9715 6071
rect 9749 6037 9783 6071
rect 9817 6037 9851 6071
rect 9886 6037 9920 6071
rect 9955 6037 9989 6071
rect 10024 6037 10058 6071
rect 10093 6037 10127 6071
rect 10162 6037 10196 6071
rect 10231 6037 10265 6071
rect 10300 6037 10334 6071
rect 10369 6037 10403 6071
rect 10438 6037 10472 6071
rect 10507 6037 10541 6071
rect 10576 6037 10610 6071
rect 10645 6037 10679 6071
rect 10714 6037 10748 6071
rect 10783 6037 10817 6071
rect 10852 6037 10886 6071
rect 10921 6037 10955 6071
rect 10990 6037 11024 6071
rect 11059 6037 11093 6071
rect 11128 6037 11162 6071
rect 11197 6037 11231 6071
rect 11266 6037 11300 6071
rect 11335 6037 11369 6071
rect 11404 6037 11438 6071
rect 11473 6037 11507 6071
rect 11542 6037 11576 6071
rect 11611 6037 11645 6071
rect 11680 6037 11714 6071
rect 11749 6037 11783 6071
rect 11818 6037 11852 6071
rect 11887 6037 11921 6071
rect 11956 6037 11990 6071
rect 12025 6037 12059 6071
rect 12094 6037 12128 6071
rect 12163 6037 12197 6071
rect 12232 6037 12266 6071
rect 12301 6037 12335 6071
rect 12370 6037 12404 6071
rect 12439 6037 12473 6071
rect 12508 6037 12542 6071
rect 12577 6037 12611 6071
rect 12646 6037 12680 6071
rect 12715 6037 12749 6071
rect 12784 6037 12818 6071
rect 12853 6037 12887 6071
rect 12922 6037 12956 6071
rect 12991 6037 13025 6071
rect 13060 6037 13094 6071
rect 13129 6037 13163 6071
rect 3373 5994 3407 6028
rect 3441 5994 3475 6028
rect 3509 5994 3543 6028
rect 3577 5994 3611 6028
rect 3645 5994 3679 6028
rect 3713 5994 3747 6028
rect 3781 5994 3815 6028
rect 3849 5994 3883 6028
rect 3917 5994 3951 6028
rect 3985 5994 4019 6028
rect 4053 5994 4087 6028
rect 4121 5994 4155 6028
rect 4189 5994 4223 6028
rect 4257 5994 4291 6028
rect 4325 5994 4359 6028
rect 4393 5994 4427 6028
rect 4461 5994 4495 6028
rect 4529 5994 4563 6028
rect 4597 5994 4631 6028
rect 4665 5994 4699 6028
rect 4733 5994 4767 6028
rect 4801 5994 4835 6028
rect 4869 5994 4903 6028
rect 4937 5994 4971 6028
rect 5005 5994 5039 6028
rect 5073 5994 5107 6028
rect 5155 5974 5189 6008
rect 5223 5974 5257 6008
rect 5291 5974 5325 6008
rect 5359 5974 5393 6008
rect 5427 5974 5461 6008
rect 5495 5974 5529 6008
rect 5563 5974 5597 6008
rect 5631 5974 5665 6008
rect 5699 5974 5733 6008
rect 5767 5974 5801 6008
rect 5835 5974 5869 6008
rect 5903 5974 5937 6008
rect 5971 5974 6005 6008
rect 6040 5977 6074 6011
rect 6108 5977 6142 6011
rect 6176 5977 6210 6011
rect 6244 5977 6278 6011
rect 6312 5977 6346 6011
rect 6380 5977 6414 6011
rect 6448 5977 6482 6011
rect 6516 5977 6550 6011
rect 6584 5977 6618 6011
rect 6652 5977 6686 6011
rect 6720 5977 6754 6011
rect 3373 5924 3407 5958
rect 3441 5924 3475 5958
rect 3509 5924 3543 5958
rect 3577 5924 3611 5958
rect 3645 5924 3679 5958
rect 3713 5924 3747 5958
rect 3781 5924 3815 5958
rect 3849 5924 3883 5958
rect 3917 5924 3951 5958
rect 3985 5924 4019 5958
rect 4053 5924 4087 5958
rect 4121 5924 4155 5958
rect 4189 5924 4223 5958
rect 4257 5924 4291 5958
rect 4325 5924 4359 5958
rect 4393 5924 4427 5958
rect 4461 5924 4495 5958
rect 4529 5924 4563 5958
rect 4597 5924 4631 5958
rect 4665 5924 4699 5958
rect 4733 5924 4767 5958
rect 4801 5924 4835 5958
rect 4869 5924 4903 5958
rect 4937 5924 4971 5958
rect 5005 5924 5039 5958
rect 5073 5924 5107 5958
rect 5155 5904 5189 5938
rect 5223 5904 5257 5938
rect 5291 5904 5325 5938
rect 5359 5904 5393 5938
rect 5427 5904 5461 5938
rect 5495 5904 5529 5938
rect 5563 5904 5597 5938
rect 5631 5904 5665 5938
rect 5699 5904 5733 5938
rect 5767 5904 5801 5938
rect 5835 5904 5869 5938
rect 5903 5904 5937 5938
rect 5971 5904 6005 5938
rect 6040 5908 6074 5942
rect 6108 5908 6142 5942
rect 6176 5908 6210 5942
rect 6244 5908 6278 5942
rect 6312 5908 6346 5942
rect 6380 5908 6414 5942
rect 6448 5908 6482 5942
rect 6516 5908 6550 5942
rect 6584 5908 6618 5942
rect 6652 5908 6686 5942
rect 6720 5908 6754 5942
rect 3373 5854 3407 5888
rect 3441 5854 3475 5888
rect 3509 5854 3543 5888
rect 3577 5854 3611 5888
rect 3645 5854 3679 5888
rect 3713 5854 3747 5888
rect 3781 5854 3815 5888
rect 3849 5854 3883 5888
rect 3917 5854 3951 5888
rect 3985 5854 4019 5888
rect 4053 5854 4087 5888
rect 4121 5854 4155 5888
rect 4189 5854 4223 5888
rect 4257 5854 4291 5888
rect 4325 5854 4359 5888
rect 4393 5854 4427 5888
rect 4461 5854 4495 5888
rect 4529 5854 4563 5888
rect 4597 5854 4631 5888
rect 4665 5854 4699 5888
rect 4733 5854 4767 5888
rect 4801 5854 4835 5888
rect 4869 5854 4903 5888
rect 4937 5854 4971 5888
rect 5005 5854 5039 5888
rect 5073 5854 5107 5888
rect 5155 5834 5189 5868
rect 5223 5834 5257 5868
rect 5291 5834 5325 5868
rect 5359 5834 5393 5868
rect 5427 5834 5461 5868
rect 5495 5834 5529 5868
rect 5563 5834 5597 5868
rect 5631 5834 5665 5868
rect 5699 5834 5733 5868
rect 5767 5834 5801 5868
rect 5835 5834 5869 5868
rect 5903 5834 5937 5868
rect 5971 5834 6005 5868
rect 6040 5839 6074 5873
rect 6108 5839 6142 5873
rect 6176 5839 6210 5873
rect 6244 5839 6278 5873
rect 6312 5839 6346 5873
rect 6380 5839 6414 5873
rect 6448 5839 6482 5873
rect 6516 5839 6550 5873
rect 6584 5839 6618 5873
rect 6652 5839 6686 5873
rect 6720 5839 6754 5873
rect 3373 5784 3407 5818
rect 3441 5784 3475 5818
rect 3509 5784 3543 5818
rect 3577 5784 3611 5818
rect 3645 5784 3679 5818
rect 3713 5784 3747 5818
rect 3781 5784 3815 5818
rect 3849 5784 3883 5818
rect 3917 5784 3951 5818
rect 3985 5784 4019 5818
rect 4053 5784 4087 5818
rect 4121 5784 4155 5818
rect 4189 5784 4223 5818
rect 4257 5784 4291 5818
rect 4325 5784 4359 5818
rect 4393 5784 4427 5818
rect 4461 5784 4495 5818
rect 4529 5784 4563 5818
rect 4597 5784 4631 5818
rect 4665 5784 4699 5818
rect 4733 5784 4767 5818
rect 4801 5784 4835 5818
rect 4869 5784 4903 5818
rect 4937 5784 4971 5818
rect 5005 5784 5039 5818
rect 5073 5784 5107 5818
rect 5155 5764 5189 5798
rect 5223 5764 5257 5798
rect 5291 5764 5325 5798
rect 5359 5764 5393 5798
rect 5427 5764 5461 5798
rect 5495 5764 5529 5798
rect 5563 5764 5597 5798
rect 5631 5764 5665 5798
rect 5699 5764 5733 5798
rect 5767 5764 5801 5798
rect 5835 5764 5869 5798
rect 5903 5764 5937 5798
rect 5971 5764 6005 5798
rect 6040 5770 6074 5804
rect 6108 5770 6142 5804
rect 6176 5770 6210 5804
rect 6244 5770 6278 5804
rect 6312 5770 6346 5804
rect 6380 5770 6414 5804
rect 6448 5770 6482 5804
rect 6516 5770 6550 5804
rect 6584 5770 6618 5804
rect 6652 5770 6686 5804
rect 6720 5770 6754 5804
rect 3373 5714 3407 5748
rect 3441 5714 3475 5748
rect 3509 5714 3543 5748
rect 3577 5714 3611 5748
rect 3645 5714 3679 5748
rect 3713 5714 3747 5748
rect 3781 5714 3815 5748
rect 3849 5714 3883 5748
rect 3917 5714 3951 5748
rect 3985 5714 4019 5748
rect 4053 5714 4087 5748
rect 4121 5714 4155 5748
rect 4189 5714 4223 5748
rect 4257 5714 4291 5748
rect 4325 5714 4359 5748
rect 4393 5714 4427 5748
rect 4461 5714 4495 5748
rect 4529 5714 4563 5748
rect 4597 5714 4631 5748
rect 4665 5714 4699 5748
rect 4733 5714 4767 5748
rect 4801 5714 4835 5748
rect 4869 5714 4903 5748
rect 4937 5714 4971 5748
rect 5005 5714 5039 5748
rect 5073 5714 5107 5748
rect 5155 5694 5189 5728
rect 5223 5694 5257 5728
rect 5291 5694 5325 5728
rect 5359 5694 5393 5728
rect 5427 5694 5461 5728
rect 5495 5694 5529 5728
rect 5563 5694 5597 5728
rect 5631 5694 5665 5728
rect 5699 5694 5733 5728
rect 5767 5694 5801 5728
rect 5835 5694 5869 5728
rect 5903 5694 5937 5728
rect 5971 5694 6005 5728
rect 6040 5701 6074 5735
rect 6108 5701 6142 5735
rect 6176 5701 6210 5735
rect 6244 5701 6278 5735
rect 6312 5701 6346 5735
rect 6380 5701 6414 5735
rect 6448 5701 6482 5735
rect 6516 5701 6550 5735
rect 6584 5701 6618 5735
rect 6652 5701 6686 5735
rect 6720 5701 6754 5735
rect 6825 5689 6859 5723
rect 6893 5689 6927 5723
rect 6961 5689 6995 5723
rect 7029 5689 7063 5723
rect 7097 5689 7131 5723
rect 7165 5689 7199 5723
rect 7233 5689 7267 5723
rect 7301 5689 7335 5723
rect 7369 5689 7403 5723
rect 7437 5689 7471 5723
rect 7505 5689 7539 5723
rect 7573 5689 7607 5723
rect 7641 5689 7675 5723
rect 7709 5689 7743 5723
rect 7777 5689 7811 5723
rect 7845 5689 7879 5723
rect 7913 5689 7947 5723
rect 7981 5689 8015 5723
rect 8049 5689 8083 5723
rect 8117 5689 8151 5723
rect 8185 5689 8219 5723
rect 8253 5689 8287 5723
rect 8321 5689 8355 5723
rect 8389 5689 8423 5723
rect 8457 5689 8491 5723
rect 8525 5689 8559 5723
rect 8593 5689 8627 5723
rect 8661 5689 8695 5723
rect 8729 5689 8763 5723
rect 8797 5689 8831 5723
rect 8865 5689 8899 5723
rect 8933 5689 8967 5723
rect 9001 5689 9035 5723
rect 9069 5689 9103 5723
rect 9137 5689 9171 5723
rect 9205 5689 9239 5723
rect 9273 5689 9307 5723
rect 9341 5689 9375 5723
rect 9409 5689 9443 5723
rect 9477 5689 9511 5723
rect 9545 5689 9579 5723
rect 9613 5689 9647 5723
rect 9681 5689 9715 5723
rect 9749 5689 9783 5723
rect 9817 5689 9851 5723
rect 9886 5689 9920 5723
rect 9955 5689 9989 5723
rect 10024 5689 10058 5723
rect 10093 5689 10127 5723
rect 10162 5689 10196 5723
rect 10231 5689 10265 5723
rect 10300 5689 10334 5723
rect 10369 5689 10403 5723
rect 10438 5689 10472 5723
rect 10507 5689 10541 5723
rect 10576 5689 10610 5723
rect 10645 5689 10679 5723
rect 10714 5689 10748 5723
rect 10783 5689 10817 5723
rect 10852 5689 10886 5723
rect 10921 5689 10955 5723
rect 10990 5689 11024 5723
rect 11059 5689 11093 5723
rect 11128 5689 11162 5723
rect 11197 5689 11231 5723
rect 11266 5689 11300 5723
rect 11335 5689 11369 5723
rect 11404 5689 11438 5723
rect 11473 5689 11507 5723
rect 11542 5689 11576 5723
rect 11611 5689 11645 5723
rect 11680 5689 11714 5723
rect 11749 5689 11783 5723
rect 11818 5689 11852 5723
rect 11887 5689 11921 5723
rect 11956 5689 11990 5723
rect 12025 5689 12059 5723
rect 12094 5689 12128 5723
rect 12163 5689 12197 5723
rect 12232 5689 12266 5723
rect 12301 5689 12335 5723
rect 12370 5689 12404 5723
rect 12439 5689 12473 5723
rect 12508 5689 12542 5723
rect 12577 5689 12611 5723
rect 12646 5689 12680 5723
rect 12715 5689 12749 5723
rect 12784 5689 12818 5723
rect 12853 5689 12887 5723
rect 12922 5689 12956 5723
rect 12991 5689 13025 5723
rect 13060 5689 13094 5723
rect 13129 5689 13163 5723
rect 3373 5644 3407 5678
rect 3441 5644 3475 5678
rect 3509 5644 3543 5678
rect 3577 5644 3611 5678
rect 3645 5644 3679 5678
rect 3713 5644 3747 5678
rect 3781 5644 3815 5678
rect 3849 5644 3883 5678
rect 3917 5644 3951 5678
rect 3985 5644 4019 5678
rect 4053 5644 4087 5678
rect 4121 5644 4155 5678
rect 4189 5644 4223 5678
rect 4257 5644 4291 5678
rect 4325 5644 4359 5678
rect 4393 5644 4427 5678
rect 4461 5644 4495 5678
rect 4529 5644 4563 5678
rect 4597 5644 4631 5678
rect 4665 5644 4699 5678
rect 4733 5644 4767 5678
rect 4801 5644 4835 5678
rect 4869 5644 4903 5678
rect 4937 5644 4971 5678
rect 5005 5644 5039 5678
rect 5073 5644 5107 5678
rect 5155 5623 5189 5657
rect 5223 5623 5257 5657
rect 5291 5623 5325 5657
rect 5359 5623 5393 5657
rect 5427 5623 5461 5657
rect 5495 5623 5529 5657
rect 5563 5623 5597 5657
rect 5631 5623 5665 5657
rect 5699 5623 5733 5657
rect 5767 5623 5801 5657
rect 5835 5623 5869 5657
rect 5903 5623 5937 5657
rect 5971 5623 6005 5657
rect 6040 5632 6074 5666
rect 6108 5632 6142 5666
rect 6176 5632 6210 5666
rect 6244 5632 6278 5666
rect 6312 5632 6346 5666
rect 6380 5632 6414 5666
rect 6448 5632 6482 5666
rect 6516 5632 6550 5666
rect 6584 5632 6618 5666
rect 6652 5632 6686 5666
rect 6720 5632 6754 5666
rect 3373 5574 3407 5608
rect 3441 5574 3475 5608
rect 3509 5574 3543 5608
rect 3577 5574 3611 5608
rect 3645 5574 3679 5608
rect 3713 5574 3747 5608
rect 3781 5574 3815 5608
rect 3849 5574 3883 5608
rect 3917 5574 3951 5608
rect 3985 5574 4019 5608
rect 4053 5574 4087 5608
rect 4121 5574 4155 5608
rect 4189 5574 4223 5608
rect 4257 5574 4291 5608
rect 4325 5574 4359 5608
rect 4393 5574 4427 5608
rect 4461 5574 4495 5608
rect 4529 5574 4563 5608
rect 4597 5574 4631 5608
rect 4665 5574 4699 5608
rect 4733 5574 4767 5608
rect 4801 5574 4835 5608
rect 4869 5574 4903 5608
rect 4937 5574 4971 5608
rect 5005 5574 5039 5608
rect 5073 5574 5107 5608
rect 5155 5552 5189 5586
rect 5223 5552 5257 5586
rect 5291 5552 5325 5586
rect 5359 5552 5393 5586
rect 5427 5552 5461 5586
rect 5495 5552 5529 5586
rect 5563 5552 5597 5586
rect 5631 5552 5665 5586
rect 5699 5552 5733 5586
rect 5767 5552 5801 5586
rect 5835 5552 5869 5586
rect 5903 5552 5937 5586
rect 5971 5552 6005 5586
rect 6040 5563 6074 5597
rect 6108 5563 6142 5597
rect 6176 5563 6210 5597
rect 6244 5563 6278 5597
rect 6312 5563 6346 5597
rect 6380 5563 6414 5597
rect 6448 5563 6482 5597
rect 6516 5563 6550 5597
rect 6584 5563 6618 5597
rect 6652 5563 6686 5597
rect 6720 5563 6754 5597
rect 3373 5504 3407 5538
rect 3441 5504 3475 5538
rect 3509 5504 3543 5538
rect 3577 5504 3611 5538
rect 3645 5504 3679 5538
rect 3713 5504 3747 5538
rect 3781 5504 3815 5538
rect 3849 5504 3883 5538
rect 3917 5504 3951 5538
rect 3985 5504 4019 5538
rect 4053 5504 4087 5538
rect 4121 5504 4155 5538
rect 4189 5504 4223 5538
rect 4257 5504 4291 5538
rect 4325 5504 4359 5538
rect 4393 5504 4427 5538
rect 4461 5504 4495 5538
rect 4529 5504 4563 5538
rect 4597 5504 4631 5538
rect 4665 5504 4699 5538
rect 4733 5504 4767 5538
rect 4801 5504 4835 5538
rect 4869 5504 4903 5538
rect 4937 5504 4971 5538
rect 5005 5504 5039 5538
rect 5073 5504 5107 5538
rect 5155 5471 5189 5505
rect 5223 5471 5257 5505
rect 5291 5471 5325 5505
rect 5359 5471 5393 5505
rect 5427 5471 5461 5505
rect 5495 5471 5529 5505
rect 5563 5471 5597 5505
rect 5631 5471 5665 5505
rect 5699 5471 5733 5505
rect 5767 5471 5801 5505
rect 5835 5471 5869 5505
rect 5903 5471 5937 5505
rect 5971 5471 6005 5505
rect 6040 5494 6074 5528
rect 6108 5494 6142 5528
rect 6176 5494 6210 5528
rect 6244 5494 6278 5528
rect 6312 5494 6346 5528
rect 6380 5494 6414 5528
rect 6448 5494 6482 5528
rect 6516 5494 6550 5528
rect 6584 5494 6618 5528
rect 6652 5494 6686 5528
rect 6720 5494 6754 5528
rect 3373 5434 3407 5468
rect 3441 5434 3475 5468
rect 3509 5434 3543 5468
rect 3577 5434 3611 5468
rect 3645 5434 3679 5468
rect 3713 5434 3747 5468
rect 3781 5434 3815 5468
rect 3849 5434 3883 5468
rect 3917 5434 3951 5468
rect 3985 5434 4019 5468
rect 4053 5434 4087 5468
rect 4121 5434 4155 5468
rect 4189 5434 4223 5468
rect 4257 5434 4291 5468
rect 4325 5434 4359 5468
rect 4393 5434 4427 5468
rect 4461 5434 4495 5468
rect 4529 5434 4563 5468
rect 4597 5434 4631 5468
rect 4665 5434 4699 5468
rect 4733 5434 4767 5468
rect 4801 5434 4835 5468
rect 4869 5434 4903 5468
rect 4937 5434 4971 5468
rect 5005 5434 5039 5468
rect 5073 5434 5107 5468
rect 3373 5364 3407 5398
rect 3441 5364 3475 5398
rect 3509 5364 3543 5398
rect 3577 5364 3611 5398
rect 3645 5364 3679 5398
rect 3713 5364 3747 5398
rect 3781 5364 3815 5398
rect 3849 5364 3883 5398
rect 3917 5364 3951 5398
rect 3985 5364 4019 5398
rect 4053 5364 4087 5398
rect 4121 5364 4155 5398
rect 4189 5364 4223 5398
rect 4257 5364 4291 5398
rect 4325 5364 4359 5398
rect 4393 5364 4427 5398
rect 4461 5364 4495 5398
rect 4529 5364 4563 5398
rect 4597 5364 4631 5398
rect 4665 5364 4699 5398
rect 4733 5364 4767 5398
rect 4801 5364 4835 5398
rect 4869 5364 4903 5398
rect 4937 5364 4971 5398
rect 5005 5364 5039 5398
rect 5073 5364 5107 5398
rect 5155 5397 5189 5431
rect 5223 5397 5257 5431
rect 5291 5397 5325 5431
rect 5359 5397 5393 5431
rect 5427 5397 5461 5431
rect 5495 5397 5529 5431
rect 5563 5397 5597 5431
rect 5631 5397 5665 5431
rect 5699 5397 5733 5431
rect 5767 5397 5801 5431
rect 5835 5397 5869 5431
rect 5903 5397 5937 5431
rect 5971 5397 6005 5431
rect 6040 5425 6074 5459
rect 6108 5425 6142 5459
rect 6176 5425 6210 5459
rect 6244 5425 6278 5459
rect 6312 5425 6346 5459
rect 6380 5425 6414 5459
rect 6448 5425 6482 5459
rect 6516 5425 6550 5459
rect 6584 5425 6618 5459
rect 6652 5425 6686 5459
rect 6720 5425 6754 5459
rect 6040 5356 6074 5390
rect 6108 5356 6142 5390
rect 6176 5356 6210 5390
rect 6244 5356 6278 5390
rect 6312 5356 6346 5390
rect 6380 5356 6414 5390
rect 6448 5356 6482 5390
rect 6516 5356 6550 5390
rect 6584 5356 6618 5390
rect 6652 5356 6686 5390
rect 6720 5356 6754 5390
rect 3373 5294 3407 5328
rect 3441 5294 3475 5328
rect 3509 5294 3543 5328
rect 3577 5294 3611 5328
rect 3645 5294 3679 5328
rect 3713 5294 3747 5328
rect 3781 5294 3815 5328
rect 3849 5294 3883 5328
rect 3917 5294 3951 5328
rect 3985 5294 4019 5328
rect 4053 5294 4087 5328
rect 4121 5294 4155 5328
rect 4189 5294 4223 5328
rect 4257 5294 4291 5328
rect 4325 5294 4359 5328
rect 4393 5294 4427 5328
rect 4461 5294 4495 5328
rect 4529 5294 4563 5328
rect 4597 5294 4631 5328
rect 4665 5294 4699 5328
rect 4733 5294 4767 5328
rect 4801 5294 4835 5328
rect 4869 5294 4903 5328
rect 4937 5294 4971 5328
rect 5005 5294 5039 5328
rect 5073 5294 5107 5328
rect 5155 5322 5189 5356
rect 5223 5322 5257 5356
rect 5291 5322 5325 5356
rect 5359 5322 5393 5356
rect 5427 5322 5461 5356
rect 5495 5322 5529 5356
rect 5563 5322 5597 5356
rect 5631 5322 5665 5356
rect 5699 5322 5733 5356
rect 5767 5322 5801 5356
rect 5835 5322 5869 5356
rect 5903 5322 5937 5356
rect 5971 5322 6005 5356
rect 6825 5341 6859 5375
rect 6893 5341 6927 5375
rect 6961 5341 6995 5375
rect 7029 5341 7063 5375
rect 7097 5341 7131 5375
rect 7165 5341 7199 5375
rect 7233 5341 7267 5375
rect 7301 5341 7335 5375
rect 7369 5341 7403 5375
rect 7437 5341 7471 5375
rect 7505 5341 7539 5375
rect 7573 5341 7607 5375
rect 7641 5341 7675 5375
rect 7709 5341 7743 5375
rect 7777 5341 7811 5375
rect 7845 5341 7879 5375
rect 7913 5341 7947 5375
rect 7981 5341 8015 5375
rect 8049 5341 8083 5375
rect 8117 5341 8151 5375
rect 8185 5341 8219 5375
rect 8253 5341 8287 5375
rect 8321 5341 8355 5375
rect 8389 5341 8423 5375
rect 8457 5341 8491 5375
rect 8525 5341 8559 5375
rect 8593 5341 8627 5375
rect 8661 5341 8695 5375
rect 8729 5341 8763 5375
rect 8797 5341 8831 5375
rect 8865 5341 8899 5375
rect 8933 5341 8967 5375
rect 9001 5341 9035 5375
rect 9069 5341 9103 5375
rect 9137 5341 9171 5375
rect 9205 5341 9239 5375
rect 9273 5341 9307 5375
rect 9341 5341 9375 5375
rect 9409 5341 9443 5375
rect 9477 5341 9511 5375
rect 9545 5341 9579 5375
rect 9613 5341 9647 5375
rect 9681 5341 9715 5375
rect 9749 5341 9783 5375
rect 9817 5341 9851 5375
rect 9886 5341 9920 5375
rect 9955 5341 9989 5375
rect 10024 5341 10058 5375
rect 10093 5341 10127 5375
rect 10162 5341 10196 5375
rect 10231 5341 10265 5375
rect 10300 5341 10334 5375
rect 10369 5341 10403 5375
rect 10438 5341 10472 5375
rect 10507 5341 10541 5375
rect 10576 5341 10610 5375
rect 10645 5341 10679 5375
rect 10714 5341 10748 5375
rect 10783 5341 10817 5375
rect 10852 5341 10886 5375
rect 10921 5341 10955 5375
rect 10990 5341 11024 5375
rect 11059 5341 11093 5375
rect 11128 5341 11162 5375
rect 11197 5341 11231 5375
rect 11266 5341 11300 5375
rect 11335 5341 11369 5375
rect 11404 5341 11438 5375
rect 11473 5341 11507 5375
rect 11542 5341 11576 5375
rect 11611 5341 11645 5375
rect 11680 5341 11714 5375
rect 11749 5341 11783 5375
rect 11818 5341 11852 5375
rect 11887 5341 11921 5375
rect 11956 5341 11990 5375
rect 12025 5341 12059 5375
rect 12094 5341 12128 5375
rect 12163 5341 12197 5375
rect 12232 5341 12266 5375
rect 12301 5341 12335 5375
rect 12370 5341 12404 5375
rect 12439 5341 12473 5375
rect 12508 5341 12542 5375
rect 12577 5341 12611 5375
rect 12646 5341 12680 5375
rect 12715 5341 12749 5375
rect 12784 5341 12818 5375
rect 12853 5341 12887 5375
rect 12922 5341 12956 5375
rect 12991 5341 13025 5375
rect 13060 5341 13094 5375
rect 13129 5341 13163 5375
rect 6040 5287 6074 5321
rect 6108 5287 6142 5321
rect 6176 5287 6210 5321
rect 6244 5287 6278 5321
rect 6312 5287 6346 5321
rect 6380 5287 6414 5321
rect 6448 5287 6482 5321
rect 6516 5287 6550 5321
rect 6584 5287 6618 5321
rect 6652 5287 6686 5321
rect 6720 5287 6754 5321
rect 3373 5223 3407 5257
rect 3441 5223 3475 5257
rect 3509 5223 3543 5257
rect 3577 5223 3611 5257
rect 3645 5223 3679 5257
rect 3713 5223 3747 5257
rect 3781 5223 3815 5257
rect 3849 5223 3883 5257
rect 3917 5223 3951 5257
rect 3985 5223 4019 5257
rect 4053 5223 4087 5257
rect 4121 5223 4155 5257
rect 4189 5223 4223 5257
rect 4257 5223 4291 5257
rect 4325 5223 4359 5257
rect 4393 5223 4427 5257
rect 4461 5223 4495 5257
rect 4529 5223 4563 5257
rect 4597 5223 4631 5257
rect 4665 5223 4699 5257
rect 4733 5223 4767 5257
rect 4801 5223 4835 5257
rect 4869 5223 4903 5257
rect 4937 5223 4971 5257
rect 5005 5223 5039 5257
rect 5073 5223 5107 5257
rect 5155 5247 5189 5281
rect 5223 5247 5257 5281
rect 5291 5247 5325 5281
rect 5359 5247 5393 5281
rect 5427 5247 5461 5281
rect 5495 5247 5529 5281
rect 5563 5247 5597 5281
rect 5631 5247 5665 5281
rect 5699 5247 5733 5281
rect 5767 5247 5801 5281
rect 5835 5247 5869 5281
rect 5903 5247 5937 5281
rect 5971 5247 6005 5281
rect 6040 5217 6074 5251
rect 6108 5217 6142 5251
rect 6176 5217 6210 5251
rect 6244 5217 6278 5251
rect 6312 5217 6346 5251
rect 6380 5217 6414 5251
rect 6448 5217 6482 5251
rect 6516 5217 6550 5251
rect 6584 5217 6618 5251
rect 6652 5217 6686 5251
rect 6720 5217 6754 5251
rect 3373 5152 3407 5186
rect 3441 5152 3475 5186
rect 3509 5152 3543 5186
rect 3577 5152 3611 5186
rect 3645 5152 3679 5186
rect 3713 5152 3747 5186
rect 3781 5152 3815 5186
rect 3849 5152 3883 5186
rect 3917 5152 3951 5186
rect 3985 5152 4019 5186
rect 4053 5152 4087 5186
rect 4121 5152 4155 5186
rect 4189 5152 4223 5186
rect 4257 5152 4291 5186
rect 4325 5152 4359 5186
rect 4393 5152 4427 5186
rect 4461 5152 4495 5186
rect 4529 5152 4563 5186
rect 4597 5152 4631 5186
rect 4665 5152 4699 5186
rect 4733 5152 4767 5186
rect 4801 5152 4835 5186
rect 4869 5152 4903 5186
rect 4937 5152 4971 5186
rect 5005 5152 5039 5186
rect 5073 5152 5107 5186
rect 5155 5172 5189 5206
rect 5223 5172 5257 5206
rect 5291 5172 5325 5206
rect 5359 5172 5393 5206
rect 5427 5172 5461 5206
rect 5495 5172 5529 5206
rect 5563 5172 5597 5206
rect 5631 5172 5665 5206
rect 5699 5172 5733 5206
rect 5767 5172 5801 5206
rect 5835 5172 5869 5206
rect 5903 5172 5937 5206
rect 5971 5172 6005 5206
rect 6040 5147 6074 5181
rect 6108 5147 6142 5181
rect 6176 5147 6210 5181
rect 6244 5147 6278 5181
rect 6312 5147 6346 5181
rect 6380 5147 6414 5181
rect 6448 5147 6482 5181
rect 6516 5147 6550 5181
rect 6584 5147 6618 5181
rect 6652 5147 6686 5181
rect 6720 5147 6754 5181
rect 3373 5081 3407 5115
rect 3441 5081 3475 5115
rect 3509 5081 3543 5115
rect 3577 5081 3611 5115
rect 3645 5081 3679 5115
rect 3713 5081 3747 5115
rect 3781 5081 3815 5115
rect 3849 5081 3883 5115
rect 3917 5081 3951 5115
rect 3985 5081 4019 5115
rect 4053 5081 4087 5115
rect 4121 5081 4155 5115
rect 4189 5081 4223 5115
rect 4257 5081 4291 5115
rect 4325 5081 4359 5115
rect 4393 5081 4427 5115
rect 4461 5081 4495 5115
rect 4529 5081 4563 5115
rect 4597 5081 4631 5115
rect 4665 5081 4699 5115
rect 4733 5081 4767 5115
rect 4801 5081 4835 5115
rect 4869 5081 4903 5115
rect 4937 5081 4971 5115
rect 5005 5081 5039 5115
rect 5073 5081 5107 5115
rect 5155 5097 5189 5131
rect 5223 5097 5257 5131
rect 5291 5097 5325 5131
rect 5359 5097 5393 5131
rect 5427 5097 5461 5131
rect 5495 5097 5529 5131
rect 5563 5097 5597 5131
rect 5631 5097 5665 5131
rect 5699 5097 5733 5131
rect 5767 5097 5801 5131
rect 5835 5097 5869 5131
rect 5903 5097 5937 5131
rect 5971 5097 6005 5131
rect 6040 5077 6074 5111
rect 6108 5077 6142 5111
rect 6176 5077 6210 5111
rect 6244 5077 6278 5111
rect 6312 5077 6346 5111
rect 6380 5077 6414 5111
rect 6448 5077 6482 5111
rect 6516 5077 6550 5111
rect 6584 5077 6618 5111
rect 6652 5077 6686 5111
rect 6720 5077 6754 5111
rect 3373 5010 3407 5044
rect 3441 5010 3475 5044
rect 3509 5010 3543 5044
rect 3577 5010 3611 5044
rect 3645 5010 3679 5044
rect 3713 5010 3747 5044
rect 3781 5010 3815 5044
rect 3849 5010 3883 5044
rect 3917 5010 3951 5044
rect 3985 5010 4019 5044
rect 4053 5010 4087 5044
rect 4121 5010 4155 5044
rect 4189 5010 4223 5044
rect 4257 5010 4291 5044
rect 4325 5010 4359 5044
rect 4393 5010 4427 5044
rect 4461 5010 4495 5044
rect 4529 5010 4563 5044
rect 4597 5010 4631 5044
rect 4665 5010 4699 5044
rect 4733 5010 4767 5044
rect 4801 5010 4835 5044
rect 4869 5010 4903 5044
rect 4937 5010 4971 5044
rect 5005 5010 5039 5044
rect 5073 5010 5107 5044
rect 5155 5022 5189 5056
rect 5223 5022 5257 5056
rect 5291 5022 5325 5056
rect 5359 5022 5393 5056
rect 5427 5022 5461 5056
rect 5495 5022 5529 5056
rect 5563 5022 5597 5056
rect 5631 5022 5665 5056
rect 5699 5022 5733 5056
rect 5767 5022 5801 5056
rect 5835 5022 5869 5056
rect 5903 5022 5937 5056
rect 5971 5022 6005 5056
rect 6040 5007 6074 5041
rect 6108 5007 6142 5041
rect 6176 5007 6210 5041
rect 6244 5007 6278 5041
rect 6312 5007 6346 5041
rect 6380 5007 6414 5041
rect 6448 5007 6482 5041
rect 6516 5007 6550 5041
rect 6584 5007 6618 5041
rect 6652 5007 6686 5041
rect 6720 5007 6754 5041
rect 3373 4939 3407 4973
rect 3441 4939 3475 4973
rect 3509 4939 3543 4973
rect 3577 4939 3611 4973
rect 3645 4939 3679 4973
rect 3713 4939 3747 4973
rect 3781 4939 3815 4973
rect 3849 4939 3883 4973
rect 3917 4939 3951 4973
rect 3985 4939 4019 4973
rect 4053 4939 4087 4973
rect 4121 4939 4155 4973
rect 4189 4939 4223 4973
rect 4257 4939 4291 4973
rect 4325 4939 4359 4973
rect 4393 4939 4427 4973
rect 4461 4939 4495 4973
rect 4529 4939 4563 4973
rect 4597 4939 4631 4973
rect 4665 4939 4699 4973
rect 4733 4939 4767 4973
rect 4801 4939 4835 4973
rect 4869 4939 4903 4973
rect 4937 4939 4971 4973
rect 5005 4939 5039 4973
rect 5073 4939 5107 4973
rect 5155 4947 5189 4981
rect 5223 4947 5257 4981
rect 5291 4947 5325 4981
rect 5359 4947 5393 4981
rect 5427 4947 5461 4981
rect 5495 4947 5529 4981
rect 5563 4947 5597 4981
rect 5631 4947 5665 4981
rect 5699 4947 5733 4981
rect 5767 4947 5801 4981
rect 5835 4947 5869 4981
rect 5903 4947 5937 4981
rect 5971 4947 6005 4981
rect 6040 4937 6074 4971
rect 6108 4937 6142 4971
rect 6176 4937 6210 4971
rect 6244 4937 6278 4971
rect 6312 4937 6346 4971
rect 6380 4937 6414 4971
rect 6448 4937 6482 4971
rect 6516 4937 6550 4971
rect 6584 4937 6618 4971
rect 6652 4937 6686 4971
rect 6720 4937 6754 4971
rect 6829 4951 6863 4985
rect 6898 4951 6932 4985
rect 6967 4951 7001 4985
rect 7036 4951 7070 4985
rect 7105 4951 7139 4985
rect 7174 4951 7208 4985
rect 7243 4951 7277 4985
rect 7312 4951 7346 4985
rect 7381 4951 7415 4985
rect 7450 4951 7484 4985
rect 7519 4951 7553 4985
rect 7588 4951 7622 4985
rect 7657 4951 7691 4985
rect 7726 4951 7760 4985
rect 7795 4951 7829 4985
rect 7864 4951 7898 4985
rect 7933 4951 7967 4985
rect 8002 4951 8036 4985
rect 8071 4951 8105 4985
rect 8140 4951 8174 4985
rect 8209 4951 8243 4985
rect 8278 4951 8312 4985
rect 8347 4951 8381 4985
rect 8416 4951 8450 4985
rect 8485 4951 8519 4985
rect 8554 4951 8588 4985
rect 3373 4868 3407 4902
rect 3441 4868 3475 4902
rect 3509 4868 3543 4902
rect 3577 4868 3611 4902
rect 3645 4868 3679 4902
rect 3713 4868 3747 4902
rect 3781 4868 3815 4902
rect 3849 4868 3883 4902
rect 3917 4868 3951 4902
rect 3985 4868 4019 4902
rect 4053 4868 4087 4902
rect 4121 4868 4155 4902
rect 4189 4868 4223 4902
rect 4257 4868 4291 4902
rect 4325 4868 4359 4902
rect 4393 4868 4427 4902
rect 4461 4868 4495 4902
rect 4529 4868 4563 4902
rect 4597 4868 4631 4902
rect 4665 4868 4699 4902
rect 4733 4868 4767 4902
rect 4801 4868 4835 4902
rect 4869 4868 4903 4902
rect 4937 4868 4971 4902
rect 5005 4868 5039 4902
rect 5073 4868 5107 4902
rect 5155 4872 5189 4906
rect 5223 4872 5257 4906
rect 5291 4872 5325 4906
rect 5359 4872 5393 4906
rect 5427 4872 5461 4906
rect 5495 4872 5529 4906
rect 5563 4872 5597 4906
rect 5631 4872 5665 4906
rect 5699 4872 5733 4906
rect 5767 4872 5801 4906
rect 5835 4872 5869 4906
rect 5903 4872 5937 4906
rect 5971 4872 6005 4906
rect 6040 4867 6074 4901
rect 6108 4867 6142 4901
rect 6176 4867 6210 4901
rect 6244 4867 6278 4901
rect 6312 4867 6346 4901
rect 6380 4867 6414 4901
rect 6448 4867 6482 4901
rect 6516 4867 6550 4901
rect 6584 4867 6618 4901
rect 6652 4867 6686 4901
rect 6720 4867 6754 4901
rect 6829 4883 6863 4917
rect 6898 4883 6932 4917
rect 6967 4883 7001 4917
rect 7036 4883 7070 4917
rect 7105 4883 7139 4917
rect 7174 4883 7208 4917
rect 7243 4883 7277 4917
rect 7312 4883 7346 4917
rect 7381 4883 7415 4917
rect 7450 4883 7484 4917
rect 7519 4883 7553 4917
rect 7588 4883 7622 4917
rect 7657 4883 7691 4917
rect 7726 4883 7760 4917
rect 7795 4883 7829 4917
rect 7864 4883 7898 4917
rect 7933 4883 7967 4917
rect 8002 4883 8036 4917
rect 8071 4883 8105 4917
rect 8140 4883 8174 4917
rect 8209 4883 8243 4917
rect 8278 4883 8312 4917
rect 8347 4883 8381 4917
rect 8416 4883 8450 4917
rect 8485 4883 8519 4917
rect 8554 4883 8588 4917
rect 3373 4797 3407 4831
rect 3441 4797 3475 4831
rect 3509 4797 3543 4831
rect 3577 4797 3611 4831
rect 3645 4797 3679 4831
rect 3713 4797 3747 4831
rect 3781 4797 3815 4831
rect 3849 4797 3883 4831
rect 3917 4797 3951 4831
rect 3985 4797 4019 4831
rect 4053 4797 4087 4831
rect 4121 4797 4155 4831
rect 4189 4797 4223 4831
rect 4257 4797 4291 4831
rect 4325 4797 4359 4831
rect 4393 4797 4427 4831
rect 4461 4797 4495 4831
rect 4529 4797 4563 4831
rect 4597 4797 4631 4831
rect 4665 4797 4699 4831
rect 4733 4797 4767 4831
rect 4801 4797 4835 4831
rect 4869 4797 4903 4831
rect 4937 4797 4971 4831
rect 5005 4797 5039 4831
rect 5073 4797 5107 4831
rect 5155 4797 5189 4831
rect 5223 4797 5257 4831
rect 5291 4797 5325 4831
rect 5359 4797 5393 4831
rect 5427 4797 5461 4831
rect 5495 4797 5529 4831
rect 5563 4797 5597 4831
rect 5631 4797 5665 4831
rect 5699 4797 5733 4831
rect 5767 4797 5801 4831
rect 5835 4797 5869 4831
rect 5903 4797 5937 4831
rect 5971 4797 6005 4831
rect 6040 4797 6074 4831
rect 6108 4797 6142 4831
rect 6176 4797 6210 4831
rect 6244 4797 6278 4831
rect 6312 4797 6346 4831
rect 6380 4797 6414 4831
rect 6448 4797 6482 4831
rect 6516 4797 6550 4831
rect 6584 4797 6618 4831
rect 6652 4797 6686 4831
rect 6720 4797 6754 4831
rect 6829 4815 6863 4849
rect 6898 4815 6932 4849
rect 6967 4815 7001 4849
rect 7036 4815 7070 4849
rect 7105 4815 7139 4849
rect 7174 4815 7208 4849
rect 7243 4815 7277 4849
rect 7312 4815 7346 4849
rect 7381 4815 7415 4849
rect 7450 4815 7484 4849
rect 7519 4815 7553 4849
rect 7588 4815 7622 4849
rect 7657 4815 7691 4849
rect 7726 4815 7760 4849
rect 7795 4815 7829 4849
rect 7864 4815 7898 4849
rect 7933 4815 7967 4849
rect 8002 4815 8036 4849
rect 8071 4815 8105 4849
rect 8140 4815 8174 4849
rect 8209 4815 8243 4849
rect 8278 4815 8312 4849
rect 8347 4815 8381 4849
rect 8416 4815 8450 4849
rect 8485 4815 8519 4849
rect 8554 4815 8588 4849
rect 8623 4815 13145 4985
rect 13197 4798 13367 6804
rect 3374 4729 3408 4763
rect 3443 4729 3477 4763
rect 3512 4729 3546 4763
rect 3581 4729 3615 4763
rect 3650 4729 3684 4763
rect 3719 4729 3753 4763
rect 3788 4729 3822 4763
rect 3857 4729 3891 4763
rect 3926 4729 3960 4763
rect 3995 4729 4029 4763
rect 4064 4729 4098 4763
rect 4133 4729 4167 4763
rect 4202 4729 4236 4763
rect 4271 4729 4305 4763
rect 4340 4729 4374 4763
rect 4409 4729 4443 4763
rect 4478 4729 4512 4763
rect 4547 4729 4581 4763
rect 4616 4729 4650 4763
rect 4685 4729 4719 4763
rect 4754 4729 4788 4763
rect 4823 4729 4857 4763
rect 4892 4729 4926 4763
rect 4961 4729 4995 4763
rect 5030 4729 5064 4763
rect 5099 4729 5133 4763
rect 5168 4729 5202 4763
rect 5237 4729 5271 4763
rect 5306 4729 5340 4763
rect 5375 4729 5409 4763
rect 5444 4729 5478 4763
rect 5513 4729 5547 4763
rect 5582 4729 5616 4763
rect 5651 4729 5685 4763
rect 5720 4729 5754 4763
rect 5789 4729 5823 4763
rect 5858 4729 5892 4763
rect 5927 4729 5961 4763
rect 5996 4729 6030 4763
rect 6065 4729 6099 4763
rect 6134 4729 6168 4763
rect 6203 4729 6237 4763
rect 6272 4729 6306 4763
rect 6341 4729 6375 4763
rect 6410 4729 6444 4763
rect 6479 4729 6513 4763
rect 6548 4729 6582 4763
rect 6617 4729 6651 4763
rect 6686 4729 6720 4763
rect 6755 4729 6789 4763
rect 6824 4729 6858 4763
rect 6893 4729 6927 4763
rect 6962 4695 10056 4763
rect 10092 4729 10126 4763
rect 10161 4729 10195 4763
rect 10230 4729 10264 4763
rect 10299 4729 10333 4763
rect 10368 4729 10402 4763
rect 10437 4729 10471 4763
rect 10506 4729 10540 4763
rect 10575 4729 10609 4763
rect 10644 4729 10678 4763
rect 10713 4729 10747 4763
rect 10782 4729 10816 4763
rect 10851 4729 10885 4763
rect 10920 4729 10954 4763
rect 10989 4729 11023 4763
rect 11058 4729 11092 4763
rect 11127 4729 11161 4763
rect 11196 4729 11230 4763
rect 11265 4729 11299 4763
rect 11334 4729 11368 4763
rect 11403 4729 11437 4763
rect 11472 4729 11506 4763
rect 11541 4729 11575 4763
rect 11610 4729 11644 4763
rect 11679 4729 11713 4763
rect 11748 4729 11782 4763
rect 11817 4729 11851 4763
rect 11886 4729 11920 4763
rect 11955 4729 11989 4763
rect 12024 4729 12058 4763
rect 12093 4729 12127 4763
rect 12162 4729 12196 4763
rect 12231 4729 12265 4763
rect 12300 4729 12334 4763
rect 12369 4729 12403 4763
rect 12438 4729 12472 4763
rect 12507 4729 12541 4763
rect 12576 4729 12610 4763
rect 12645 4729 12679 4763
rect 12714 4729 12748 4763
rect 12783 4729 12817 4763
rect 12852 4729 12886 4763
rect 12921 4729 12955 4763
rect 12990 4729 13024 4763
rect 13059 4729 13093 4763
rect 13128 4729 13162 4763
rect 13197 4729 13231 4763
rect 13265 4730 13367 4798
rect 13333 4696 13367 4730
rect 3408 4661 3442 4695
rect 3477 4661 3511 4695
rect 3546 4661 3580 4695
rect 3615 4661 3649 4695
rect 3684 4661 3718 4695
rect 3753 4661 3787 4695
rect 3822 4661 3856 4695
rect 3891 4661 3925 4695
rect 3960 4661 3994 4695
rect 4029 4661 4063 4695
rect 4098 4661 4132 4695
rect 4167 4661 4201 4695
rect 4236 4661 4270 4695
rect 4305 4661 4339 4695
rect 4374 4661 4408 4695
rect 4443 4661 4477 4695
rect 4512 4661 4546 4695
rect 4581 4661 4615 4695
rect 4650 4661 4684 4695
rect 3340 4623 3374 4657
rect 3408 4588 3442 4622
rect 3476 4593 3510 4627
rect 3545 4593 3579 4627
rect 3614 4593 3648 4627
rect 3683 4593 3717 4627
rect 3752 4593 3786 4627
rect 3821 4593 3855 4627
rect 3890 4593 3924 4627
rect 3959 4593 3993 4627
rect 4028 4593 4062 4627
rect 4097 4593 4131 4627
rect 4166 4593 4200 4627
rect 4235 4593 4269 4627
rect 4304 4593 4338 4627
rect 4373 4593 4407 4627
rect 4442 4593 4476 4627
rect 4511 4593 4545 4627
rect 4580 4593 4614 4627
rect 4649 4593 4683 4627
rect 4718 4593 10056 4695
rect 10091 4661 10125 4695
rect 10160 4661 10194 4695
rect 10229 4661 10263 4695
rect 10298 4661 10332 4695
rect 10367 4661 10401 4695
rect 10436 4661 10470 4695
rect 10505 4661 10539 4695
rect 10574 4661 10608 4695
rect 10643 4661 10677 4695
rect 10712 4661 10746 4695
rect 10781 4661 10815 4695
rect 10850 4661 10884 4695
rect 10919 4661 10953 4695
rect 10988 4661 11022 4695
rect 11057 4661 11091 4695
rect 11126 4661 11160 4695
rect 11195 4661 11229 4695
rect 11264 4661 11298 4695
rect 11333 4661 11367 4695
rect 11402 4661 11436 4695
rect 11471 4661 11505 4695
rect 11540 4661 11574 4695
rect 11609 4661 11643 4695
rect 11678 4661 11712 4695
rect 11747 4661 11781 4695
rect 11816 4661 11850 4695
rect 11885 4661 11919 4695
rect 11954 4661 11988 4695
rect 12023 4661 12057 4695
rect 12092 4661 12126 4695
rect 12161 4661 12195 4695
rect 12230 4661 12264 4695
rect 12299 4661 12333 4695
rect 12368 4661 12402 4695
rect 12437 4661 12471 4695
rect 12506 4661 12540 4695
rect 12575 4661 12609 4695
rect 12644 4661 12678 4695
rect 12713 4661 12747 4695
rect 12782 4661 12816 4695
rect 12851 4661 12885 4695
rect 12920 4661 12954 4695
rect 12989 4661 13023 4695
rect 13058 4661 13092 4695
rect 13127 4661 13161 4695
rect 13196 4661 13230 4695
rect 13265 4661 13299 4695
rect 13333 4627 13367 4661
rect 10091 4593 10125 4627
rect 10160 4593 10194 4627
rect 10229 4593 10263 4627
rect 10298 4593 10332 4627
rect 10367 4593 10401 4627
rect 10436 4593 10470 4627
rect 10505 4593 10539 4627
rect 10574 4593 10608 4627
rect 10643 4593 10677 4627
rect 10712 4593 10746 4627
rect 10781 4593 10815 4627
rect 10850 4593 10884 4627
rect 10919 4593 10953 4627
rect 10987 4593 11021 4627
rect 11055 4593 11089 4627
rect 11123 4593 11157 4627
rect 11191 4593 11225 4627
rect 11259 4593 11293 4627
rect 11327 4593 11361 4627
rect 11395 4593 11429 4627
rect 11463 4593 11497 4627
rect 11531 4593 11565 4627
rect 11599 4593 11633 4627
rect 11667 4593 11701 4627
rect 11735 4593 11769 4627
rect 11803 4593 11837 4627
rect 11871 4593 11905 4627
rect 11939 4593 11973 4627
rect 12007 4593 12041 4627
rect 12075 4593 12109 4627
rect 12143 4593 12177 4627
rect 12211 4593 12245 4627
rect 12279 4593 12313 4627
rect 12347 4593 12381 4627
rect 12415 4593 12449 4627
rect 12483 4593 12517 4627
rect 12551 4593 12585 4627
rect 12619 4593 12653 4627
rect 12687 4593 12721 4627
rect 12755 4593 12789 4627
rect 12823 4593 12857 4627
rect 12891 4593 12925 4627
rect 12959 4593 12993 4627
rect 13027 4593 13061 4627
rect 13095 4593 13129 4627
rect 13163 4593 13197 4627
rect 13231 4593 13265 4627
rect 3340 4553 3374 4587
rect 3340 4483 3374 4517
rect 3408 4515 3442 4549
rect 3476 4523 3510 4557
rect 3340 4413 3374 4447
rect 3408 4442 3442 4476
rect 3476 4453 3510 4487
rect 3340 4343 3374 4377
rect 3408 4369 3442 4403
rect 3476 4383 3510 4417
rect 3340 4273 3374 4307
rect 3408 4296 3442 4330
rect 3476 4313 3510 4347
rect 3340 4203 3374 4237
rect 3408 4222 3442 4256
rect 3476 4243 3510 4277
rect 3340 4133 3374 4167
rect 3408 4148 3442 4182
rect 3476 4173 3510 4207
rect 3340 4062 3374 4096
rect 3408 4074 3442 4108
rect 3476 4102 3510 4136
rect 3340 3991 3374 4025
rect 3408 4000 3442 4034
rect 3476 4031 3510 4065
rect 3476 3960 3510 3994
rect -1 3920 33 3954
rect 68 3920 102 3954
rect 137 3920 171 3954
rect 206 3920 240 3954
rect 275 3920 309 3954
rect 344 3920 378 3954
rect 413 3920 447 3954
rect 482 3920 516 3954
rect 551 3920 585 3954
rect 620 3886 3374 3954
rect 3408 3926 3442 3960
rect 3476 3889 3510 3923
rect -1 3852 33 3886
rect 68 3852 102 3886
rect 137 3852 171 3886
rect 206 3852 240 3886
rect 275 3852 309 3886
rect 344 3852 378 3886
rect 413 3852 447 3886
rect 482 3852 516 3886
rect 551 3852 585 3886
rect 620 3852 3442 3886
rect -1 3784 33 3818
rect 68 3784 102 3818
rect 137 3784 171 3818
rect 206 3784 240 3818
rect 275 3784 309 3818
rect 344 3784 378 3818
rect 413 3784 447 3818
rect 482 3784 516 3818
rect 551 3784 585 3818
rect 620 3784 654 3818
rect 689 3784 723 3818
rect 758 3784 792 3818
rect 827 3784 861 3818
rect 896 3784 930 3818
rect 965 3784 999 3818
rect 1034 3784 1068 3818
rect 1103 3784 1137 3818
rect 1172 3784 1206 3818
rect 1241 3784 1275 3818
rect 1310 3784 1344 3818
rect 1379 3784 1413 3818
rect 1448 3784 1482 3818
rect 1517 3784 1551 3818
rect 1586 3784 1620 3818
rect 1655 3784 1689 3818
rect 1724 3784 1758 3818
rect 1793 3784 1827 3818
rect 1862 3784 1896 3818
rect 1931 3784 1965 3818
rect 2000 3784 2034 3818
rect 2069 3784 2103 3818
rect 2138 3784 2172 3818
rect 2207 3784 2241 3818
rect 2276 3784 2310 3818
rect 2345 3784 2379 3818
rect 2414 3784 2448 3818
rect 2483 3784 2517 3818
rect 2552 3784 2586 3818
rect 2621 3784 2655 3818
rect 2690 3784 2724 3818
rect 2759 3784 2793 3818
rect 2828 3784 2862 3818
rect 2897 3784 2931 3818
rect 2966 3784 3408 3852
rect 3476 3818 3510 3852
rect 19091 2213 19125 2247
rect 19159 2213 19193 2247
rect 19091 2142 19125 2176
rect 19159 2142 19193 2176
rect 19091 2071 19125 2105
rect 19159 2071 19193 2105
rect 19091 2000 19125 2034
rect 19159 2000 19193 2034
rect 19091 1929 19125 1963
rect 19159 1929 19193 1963
rect 19091 1858 19125 1892
rect 19159 1858 19193 1892
rect 19091 1787 19125 1821
rect 19159 1787 19193 1821
rect 19091 1716 19125 1750
rect 19159 1716 19193 1750
rect 19091 1645 19125 1679
rect 19159 1645 19193 1679
rect 19091 1574 19125 1608
rect 19159 1574 19193 1608
rect 19091 1503 19125 1537
rect 19159 1503 19193 1537
rect 19091 1432 19125 1466
rect 19159 1432 19193 1466
rect 19091 1362 19125 1396
rect 19159 1362 19193 1396
rect 19091 1292 19125 1326
rect 19159 1292 19193 1326
rect 19091 1222 19125 1256
rect 19159 1222 19193 1256
rect 19091 1152 19125 1186
rect 19159 1152 19193 1186
rect 19091 1082 19125 1116
rect 19159 1082 19193 1116
rect 19091 1012 19125 1046
rect 19159 1012 19193 1046
rect 19091 942 19125 976
rect 19159 942 19193 976
<< poly >>
rect 5776 6606 5891 6622
rect 5776 6572 5792 6606
rect 5826 6572 5891 6606
rect 5776 6538 5891 6572
rect 5776 6504 5792 6538
rect 5826 6504 5891 6538
rect 5776 6470 5891 6504
rect 5776 6436 5792 6470
rect 5826 6436 5891 6470
rect 5776 6422 5891 6436
rect 6457 6606 6572 6622
rect 6457 6572 6522 6606
rect 6556 6572 6572 6606
rect 6457 6538 6572 6572
rect 6457 6504 6522 6538
rect 6556 6504 6572 6538
rect 6457 6470 6572 6504
rect 6457 6436 6522 6470
rect 6556 6436 6572 6470
rect 6457 6422 6572 6436
rect 5776 6420 5842 6422
rect 6506 6420 6572 6422
rect 6836 6279 6902 6295
rect 6836 6245 6852 6279
rect 6886 6278 6902 6279
rect 13109 6279 13175 6295
rect 13109 6278 13125 6279
rect 6886 6245 6911 6278
rect 6836 6211 6911 6245
rect 6836 6177 6852 6211
rect 6886 6178 6911 6211
rect 13100 6245 13125 6278
rect 13159 6245 13175 6279
rect 13100 6211 13175 6245
rect 13100 6178 13125 6211
rect 6886 6177 6902 6178
rect 6836 6161 6902 6177
rect 13109 6177 13125 6178
rect 13159 6177 13175 6211
rect 13109 6161 13175 6177
rect 6836 5930 6902 5946
rect 13109 5931 13175 5947
rect 13109 5930 13125 5931
rect 6836 5896 6852 5930
rect 6886 5896 6911 5930
rect 6836 5862 6911 5896
rect 6836 5828 6852 5862
rect 6886 5830 6911 5862
rect 13100 5897 13125 5930
rect 13159 5897 13175 5931
rect 13100 5863 13175 5897
rect 13100 5830 13125 5863
rect 6886 5828 6902 5830
rect 6836 5812 6902 5828
rect 13109 5829 13125 5830
rect 13159 5829 13175 5863
rect 13109 5813 13175 5829
rect 6836 5583 6902 5599
rect 6836 5549 6852 5583
rect 6886 5582 6902 5583
rect 13109 5583 13175 5599
rect 13109 5582 13125 5583
rect 6886 5549 6911 5582
rect 6836 5515 6911 5549
rect 6836 5481 6852 5515
rect 6886 5482 6911 5515
rect 13100 5549 13125 5582
rect 13159 5549 13175 5583
rect 13100 5515 13175 5549
rect 13100 5482 13125 5515
rect 6886 5481 6902 5482
rect 6836 5465 6902 5481
rect 13109 5481 13125 5482
rect 13159 5481 13175 5515
rect 13109 5465 13175 5481
rect 6836 5235 6902 5251
rect 6836 5201 6852 5235
rect 6886 5234 6902 5235
rect 13109 5235 13175 5251
rect 13109 5234 13125 5235
rect 6886 5201 6911 5234
rect 6836 5167 6911 5201
rect 6836 5133 6852 5167
rect 6886 5134 6911 5167
rect 13100 5201 13125 5234
rect 13159 5201 13175 5235
rect 13100 5167 13175 5201
rect 13100 5134 13125 5167
rect 6886 5133 6902 5134
rect 6836 5117 6902 5133
rect 13109 5133 13125 5134
rect 13159 5133 13175 5167
rect 13109 5117 13175 5133
<< polycont >>
rect 5792 6572 5826 6606
rect 5792 6504 5826 6538
rect 5792 6436 5826 6470
rect 6522 6572 6556 6606
rect 6522 6504 6556 6538
rect 6522 6436 6556 6470
rect 6852 6245 6886 6279
rect 6852 6177 6886 6211
rect 13125 6245 13159 6279
rect 13125 6177 13159 6211
rect 6852 5896 6886 5930
rect 6852 5828 6886 5862
rect 13125 5897 13159 5931
rect 13125 5829 13159 5863
rect 6852 5549 6886 5583
rect 6852 5481 6886 5515
rect 13125 5549 13159 5583
rect 13125 5481 13159 5515
rect 6852 5201 6886 5235
rect 6852 5133 6886 5167
rect 13125 5201 13159 5235
rect 13125 5133 13159 5167
<< locali >>
rect -25 6906 -1 6940
rect 33 6906 68 6940
rect 102 6906 137 6940
rect 171 6906 206 6940
rect 240 6906 275 6940
rect 309 6906 344 6940
rect 378 6906 413 6940
rect 447 6906 482 6940
rect 516 6906 551 6940
rect 585 6906 620 6940
rect 654 6906 689 6940
rect 723 6906 758 6940
rect 792 6906 827 6940
rect 861 6908 896 6940
rect 930 6908 965 6940
rect 999 6908 1034 6940
rect 1068 6908 1103 6940
rect 1137 6908 1172 6940
rect 1206 6908 1241 6940
rect 1275 6908 1310 6940
rect 1344 6908 1379 6940
rect 861 6906 865 6908
rect 930 6906 938 6908
rect 999 6906 1011 6908
rect 1068 6906 1084 6908
rect 1137 6906 1157 6908
rect 1206 6906 1230 6908
rect 1275 6906 1303 6908
rect 1344 6906 1376 6908
rect 1413 6906 1448 6940
rect 1482 6908 1517 6940
rect 1551 6908 1586 6940
rect 1620 6908 1655 6940
rect 1689 6908 1724 6940
rect 1758 6908 1793 6940
rect 1827 6908 1862 6940
rect 10056 6908 10090 6940
rect 10124 6908 10158 6940
rect 10192 6908 10226 6940
rect 10260 6908 10294 6940
rect 10328 6908 10362 6940
rect 10396 6908 10430 6940
rect 10464 6908 10498 6940
rect 10532 6908 10566 6940
rect 10600 6908 10634 6940
rect 10668 6908 10702 6940
rect 10736 6908 10770 6940
rect 10804 6908 10838 6940
rect 10872 6908 10906 6940
rect 10940 6908 10974 6940
rect 11008 6908 11042 6940
rect 11076 6908 11110 6940
rect 11144 6908 11178 6940
rect 11212 6908 11246 6940
rect 11280 6908 11314 6940
rect 11348 6908 11382 6940
rect 11416 6908 11450 6940
rect 11484 6908 11518 6940
rect 11552 6908 11586 6940
rect 11620 6908 11654 6940
rect 11688 6908 11722 6940
rect 11756 6908 11790 6940
rect 11824 6908 11858 6940
rect 11892 6908 11926 6940
rect 11960 6908 11994 6940
rect 12028 6908 12062 6940
rect 12096 6908 12130 6940
rect 12164 6908 12198 6940
rect 12232 6908 12266 6940
rect 12300 6908 12334 6940
rect 12368 6908 12402 6940
rect 12436 6908 12471 6940
rect 12505 6908 12540 6940
rect 12574 6908 12609 6940
rect 12643 6908 12678 6940
rect 12712 6908 12747 6940
rect 12781 6908 12816 6940
rect 12850 6908 12885 6940
rect 12919 6908 12954 6940
rect 12988 6908 13023 6940
rect 13057 6908 13092 6940
rect 13126 6908 13161 6940
rect 13195 6908 13230 6940
rect 13264 6908 13299 6940
rect 1483 6906 1517 6908
rect 1556 6906 1586 6908
rect 1629 6906 1655 6908
rect 1702 6906 1724 6908
rect 1775 6906 1793 6908
rect -25 6874 865 6906
rect 899 6874 938 6906
rect 972 6874 1011 6906
rect 1045 6874 1084 6906
rect 1118 6874 1157 6906
rect 1191 6874 1230 6906
rect 1264 6874 1303 6906
rect 1337 6874 1376 6906
rect 1410 6874 1449 6906
rect 1483 6874 1522 6906
rect 1556 6874 1595 6906
rect 1629 6874 1668 6906
rect 1702 6874 1741 6906
rect 1775 6874 1814 6906
rect 1848 6874 1862 6908
rect -25 6872 1862 6874
rect -25 6838 -1 6872
rect 33 6838 68 6872
rect 102 6838 137 6872
rect 171 6838 206 6872
rect 240 6838 275 6872
rect 309 6838 344 6872
rect 378 6838 413 6872
rect 447 6838 482 6872
rect 516 6838 551 6872
rect 585 6838 620 6872
rect 654 6838 689 6872
rect 723 6838 758 6872
rect 792 6838 827 6872
rect 861 6838 896 6872
rect 930 6838 965 6872
rect 999 6838 1034 6872
rect 1068 6838 1103 6872
rect 1137 6838 1172 6872
rect 1206 6838 1241 6872
rect 1275 6838 1310 6872
rect 1344 6838 1379 6872
rect 1413 6838 1448 6872
rect 1482 6838 1517 6872
rect 1551 6838 1586 6872
rect 1620 6838 1655 6872
rect 1689 6838 1724 6872
rect 1758 6838 1793 6872
rect 1827 6838 1862 6872
rect -25 6836 1862 6838
rect -25 6804 865 6836
rect 899 6804 938 6836
rect 972 6804 1011 6836
rect 1045 6804 1084 6836
rect 1118 6804 1157 6836
rect 1191 6804 1230 6836
rect 1264 6804 1303 6836
rect 1337 6804 1376 6836
rect 1410 6804 1449 6836
rect 1483 6804 1522 6836
rect 1556 6804 1595 6836
rect 1629 6804 1668 6836
rect 1702 6804 1741 6836
rect 1775 6804 1814 6836
rect -25 6770 -1 6804
rect 33 6770 68 6804
rect 102 6770 137 6804
rect 171 6770 206 6804
rect 240 6770 275 6804
rect 309 6770 344 6804
rect 378 6770 413 6804
rect 447 6770 482 6804
rect 516 6770 551 6804
rect 585 6770 620 6804
rect 654 6770 689 6804
rect 723 6770 758 6804
rect 792 6770 827 6804
rect 861 6802 865 6804
rect 930 6802 938 6804
rect 999 6802 1011 6804
rect 1068 6802 1084 6804
rect 1137 6802 1157 6804
rect 1206 6802 1230 6804
rect 1275 6802 1303 6804
rect 1344 6802 1376 6804
rect 861 6770 896 6802
rect 930 6770 965 6802
rect 999 6770 1034 6802
rect 1068 6770 1103 6802
rect 1137 6770 1172 6802
rect 1206 6770 1241 6802
rect 1275 6770 1310 6802
rect 1344 6770 1379 6802
rect 1413 6770 1448 6804
rect 1483 6802 1517 6804
rect 1556 6802 1586 6804
rect 1629 6802 1655 6804
rect 1702 6802 1724 6804
rect 1775 6802 1793 6804
rect 1848 6802 1862 6836
rect 13333 6906 13367 6940
rect 13302 6838 13367 6906
rect 1482 6770 1517 6802
rect 1551 6770 1586 6802
rect 1620 6770 1655 6802
rect 1689 6770 1724 6802
rect 1758 6770 1793 6802
rect 1827 6770 1862 6802
rect 10056 6770 10091 6802
rect 10125 6770 10160 6802
rect 10194 6770 10229 6802
rect 10263 6770 10298 6802
rect 10332 6770 10367 6802
rect 10401 6770 10436 6802
rect 10470 6770 10505 6802
rect 10539 6770 10574 6802
rect 10608 6770 10643 6802
rect 10677 6770 10712 6802
rect 10746 6770 10781 6802
rect 10815 6770 10850 6802
rect 10884 6770 10919 6802
rect 10953 6770 10988 6802
rect 11022 6770 11057 6802
rect 11091 6770 11126 6802
rect 11160 6770 11195 6802
rect 11229 6770 11264 6802
rect 11298 6770 11333 6802
rect 11367 6770 11402 6802
rect 11436 6770 11471 6802
rect 11505 6770 11540 6802
rect 11574 6770 11609 6802
rect 11643 6770 11678 6802
rect 11712 6770 11747 6802
rect 11781 6770 11816 6802
rect 11850 6770 11885 6802
rect 11919 6770 11954 6802
rect 11988 6770 12023 6802
rect 12057 6770 12092 6802
rect 12126 6770 12161 6802
rect 12195 6770 12230 6802
rect 12264 6770 12299 6802
rect 12333 6770 12368 6802
rect 12402 6770 12437 6802
rect 12471 6770 12506 6802
rect 12540 6770 12575 6802
rect 12609 6770 12644 6802
rect 12678 6770 12713 6802
rect 12747 6770 12782 6802
rect 12816 6770 12851 6802
rect 12885 6770 12920 6802
rect 12954 6770 12989 6802
rect 13023 6770 13058 6802
rect 13092 6770 13127 6802
rect 13161 6770 13197 6802
rect 2533 6751 13197 6770
rect 3340 6728 5584 6751
rect 3340 6694 3373 6728
rect 3407 6694 3441 6728
rect 3475 6694 3509 6728
rect 3543 6694 3577 6728
rect 3611 6694 3645 6728
rect 3679 6694 3713 6728
rect 3747 6694 3781 6728
rect 3815 6694 3849 6728
rect 3883 6694 3917 6728
rect 3951 6694 3985 6728
rect 4019 6694 4053 6728
rect 4087 6694 4121 6728
rect 4155 6694 4189 6728
rect 4223 6694 4257 6728
rect 4291 6694 4325 6728
rect 4359 6694 4393 6728
rect 4427 6694 4461 6728
rect 4495 6694 4529 6728
rect 4563 6694 4597 6728
rect 4631 6694 4665 6728
rect 4699 6694 4733 6728
rect 4767 6694 4801 6728
rect 4835 6694 4869 6728
rect 4903 6694 4937 6728
rect 4971 6694 5005 6728
rect 5039 6694 5073 6728
rect 5107 6695 5584 6728
rect 5107 6694 5180 6695
rect 3340 6661 5180 6694
rect 5214 6661 5248 6695
rect 5282 6661 5316 6695
rect 5350 6661 5384 6695
rect 5418 6661 5452 6695
rect 5486 6661 5520 6695
rect 5554 6661 5584 6695
rect 3340 6658 5584 6661
rect 3340 6624 3373 6658
rect 3407 6624 3441 6658
rect 3475 6624 3509 6658
rect 3543 6624 3577 6658
rect 3611 6624 3645 6658
rect 3679 6624 3713 6658
rect 3747 6624 3781 6658
rect 3815 6624 3849 6658
rect 3883 6624 3917 6658
rect 3951 6624 3985 6658
rect 4019 6624 4053 6658
rect 4087 6624 4121 6658
rect 4155 6624 4189 6658
rect 4223 6624 4257 6658
rect 4291 6624 4325 6658
rect 4359 6624 4393 6658
rect 4427 6624 4461 6658
rect 4495 6624 4529 6658
rect 4563 6624 4597 6658
rect 4631 6624 4665 6658
rect 4699 6624 4733 6658
rect 4767 6624 4801 6658
rect 4835 6624 4869 6658
rect 4903 6624 4937 6658
rect 4971 6624 5005 6658
rect 5039 6624 5073 6658
rect 5107 6625 5584 6658
rect 5870 6667 6412 6751
rect 6781 6736 6815 6751
rect 5904 6633 5945 6667
rect 5979 6633 6020 6667
rect 6054 6633 6095 6667
rect 6129 6633 6170 6667
rect 6204 6633 6245 6667
rect 6279 6633 6319 6667
rect 6353 6633 6393 6667
rect 6781 6663 6815 6702
rect 5107 6624 5180 6625
rect 3340 6591 5180 6624
rect 5214 6591 5248 6625
rect 5282 6591 5316 6625
rect 5350 6591 5384 6625
rect 5418 6591 5452 6625
rect 5486 6591 5520 6625
rect 5554 6591 5584 6625
rect 6522 6606 6556 6622
rect 3340 6588 5584 6591
rect 3340 6554 3373 6588
rect 3407 6554 3441 6588
rect 3475 6554 3509 6588
rect 3543 6554 3577 6588
rect 3611 6554 3645 6588
rect 3679 6554 3713 6588
rect 3747 6554 3781 6588
rect 3815 6554 3849 6588
rect 3883 6554 3917 6588
rect 3951 6554 3985 6588
rect 4019 6554 4053 6588
rect 4087 6554 4121 6588
rect 4155 6554 4189 6588
rect 4223 6554 4257 6588
rect 4291 6554 4325 6588
rect 4359 6554 4393 6588
rect 4427 6554 4461 6588
rect 4495 6554 4529 6588
rect 4563 6554 4597 6588
rect 4631 6554 4665 6588
rect 4699 6554 4733 6588
rect 4767 6554 4801 6588
rect 4835 6554 4869 6588
rect 4903 6554 4937 6588
rect 4971 6554 5005 6588
rect 5039 6554 5073 6588
rect 5107 6556 5584 6588
rect 5107 6554 5180 6556
rect 3340 6522 5180 6554
rect 5214 6522 5248 6556
rect 5282 6522 5316 6556
rect 5350 6522 5384 6556
rect 5418 6522 5452 6556
rect 5486 6522 5520 6556
rect 5554 6522 5584 6556
rect 3340 6518 5584 6522
rect 3340 6484 3373 6518
rect 3407 6484 3441 6518
rect 3475 6484 3509 6518
rect 3543 6484 3577 6518
rect 3611 6484 3645 6518
rect 3679 6484 3713 6518
rect 3747 6484 3781 6518
rect 3815 6484 3849 6518
rect 3883 6484 3917 6518
rect 3951 6484 3985 6518
rect 4019 6484 4053 6518
rect 4087 6484 4121 6518
rect 4155 6484 4189 6518
rect 4223 6484 4257 6518
rect 4291 6484 4325 6518
rect 4359 6484 4393 6518
rect 4427 6484 4461 6518
rect 4495 6484 4529 6518
rect 4563 6484 4597 6518
rect 4631 6484 4665 6518
rect 4699 6484 4733 6518
rect 4767 6484 4801 6518
rect 4835 6484 4869 6518
rect 4903 6484 4937 6518
rect 4971 6484 5005 6518
rect 5039 6484 5073 6518
rect 5107 6487 5584 6518
rect 5107 6484 5180 6487
rect 3340 6453 5180 6484
rect 5214 6453 5248 6487
rect 5282 6453 5316 6487
rect 5350 6453 5384 6487
rect 5418 6453 5452 6487
rect 5486 6453 5520 6487
rect 5554 6453 5584 6487
rect 3340 6448 5584 6453
rect 3340 6414 3373 6448
rect 3407 6414 3441 6448
rect 3475 6414 3509 6448
rect 3543 6414 3577 6448
rect 3611 6414 3645 6448
rect 3679 6414 3713 6448
rect 3747 6414 3781 6448
rect 3815 6414 3849 6448
rect 3883 6414 3917 6448
rect 3951 6414 3985 6448
rect 4019 6414 4053 6448
rect 4087 6414 4121 6448
rect 4155 6414 4189 6448
rect 4223 6414 4257 6448
rect 4291 6414 4325 6448
rect 4359 6414 4393 6448
rect 4427 6414 4461 6448
rect 4495 6414 4529 6448
rect 4563 6414 4597 6448
rect 4631 6414 4665 6448
rect 4699 6414 4733 6448
rect 4767 6414 4801 6448
rect 4835 6414 4869 6448
rect 4903 6414 4937 6448
rect 4971 6414 5005 6448
rect 5039 6414 5073 6448
rect 5107 6418 5584 6448
rect 5776 6572 5792 6606
rect 5826 6599 5842 6606
rect 5826 6572 6522 6599
rect 5776 6563 6556 6572
rect 5776 6504 5792 6563
rect 5826 6504 6522 6563
rect 5776 6491 6556 6504
rect 5776 6436 5792 6491
rect 5826 6445 6522 6491
rect 5826 6436 5842 6445
rect 6522 6420 6556 6436
rect 6781 6591 6815 6629
rect 6781 6519 6815 6557
rect 6781 6448 6815 6485
rect 9283 6720 13197 6751
rect 9283 6448 9317 6720
rect 13159 6482 13197 6720
rect 5107 6414 5180 6418
rect 3340 6384 5180 6414
rect 5214 6384 5248 6418
rect 5282 6384 5316 6418
rect 5350 6384 5384 6418
rect 5418 6384 5452 6418
rect 5486 6384 5520 6418
rect 5554 6384 5584 6418
rect 6781 6414 6825 6448
rect 6859 6414 6893 6448
rect 6927 6414 6961 6448
rect 6995 6414 7029 6448
rect 7063 6414 7097 6448
rect 7131 6414 7165 6448
rect 7199 6414 7233 6448
rect 7267 6414 7301 6448
rect 7335 6414 7369 6448
rect 7403 6414 7437 6448
rect 7471 6414 7505 6448
rect 7539 6414 7573 6448
rect 7607 6414 7641 6448
rect 7675 6414 7709 6448
rect 7743 6414 7777 6448
rect 7811 6414 7845 6448
rect 7879 6414 7913 6448
rect 7947 6414 7981 6448
rect 8015 6414 8049 6448
rect 8083 6414 8117 6448
rect 8151 6414 8185 6448
rect 8219 6414 8253 6448
rect 8287 6414 8321 6448
rect 8355 6414 8389 6448
rect 8423 6414 8457 6448
rect 8491 6414 8525 6448
rect 8559 6414 8593 6448
rect 8627 6414 8661 6448
rect 8695 6414 8729 6448
rect 8763 6414 8797 6448
rect 8831 6414 8865 6448
rect 8899 6414 8933 6448
rect 8967 6414 9001 6448
rect 9035 6414 9069 6448
rect 9103 6414 9137 6448
rect 9171 6414 9205 6448
rect 9239 6414 9273 6448
rect 9307 6414 9317 6448
rect 9851 6448 13197 6482
rect 9851 6414 9886 6448
rect 9920 6414 9955 6448
rect 9989 6414 10024 6448
rect 10058 6414 10093 6448
rect 10127 6414 10162 6448
rect 10196 6414 10231 6448
rect 10265 6414 10300 6448
rect 10334 6414 10369 6448
rect 10403 6414 10438 6448
rect 10472 6414 10507 6448
rect 10541 6414 10576 6448
rect 10610 6414 10645 6448
rect 10679 6414 10714 6448
rect 10748 6414 10783 6448
rect 10817 6414 10852 6448
rect 10886 6414 10921 6448
rect 10955 6414 10990 6448
rect 11024 6414 11059 6448
rect 11093 6414 11128 6448
rect 11162 6414 11197 6448
rect 11231 6414 11266 6448
rect 11300 6414 11335 6448
rect 11369 6414 11404 6448
rect 11438 6414 11473 6448
rect 11507 6414 11542 6448
rect 11576 6414 11611 6448
rect 11645 6414 11680 6448
rect 11714 6414 11749 6448
rect 11783 6414 11818 6448
rect 11852 6414 11887 6448
rect 11921 6414 11956 6448
rect 11990 6414 12025 6448
rect 12059 6414 12094 6448
rect 12128 6414 12163 6448
rect 12197 6414 12232 6448
rect 12266 6414 12301 6448
rect 12335 6414 12370 6448
rect 12404 6414 12439 6448
rect 12473 6414 12508 6448
rect 12542 6414 12577 6448
rect 12611 6414 12646 6448
rect 12680 6414 12715 6448
rect 12749 6414 12784 6448
rect 12818 6414 12853 6448
rect 12887 6414 12922 6448
rect 12956 6414 12991 6448
rect 13025 6414 13060 6448
rect 13094 6414 13129 6448
rect 13163 6414 13197 6448
rect 3340 6378 5584 6384
rect 3340 6344 3373 6378
rect 3407 6344 3441 6378
rect 3475 6344 3509 6378
rect 3543 6344 3577 6378
rect 3611 6344 3645 6378
rect 3679 6344 3713 6378
rect 3747 6344 3781 6378
rect 3815 6344 3849 6378
rect 3883 6344 3917 6378
rect 3951 6344 3985 6378
rect 4019 6344 4053 6378
rect 4087 6344 4121 6378
rect 4155 6344 4189 6378
rect 4223 6344 4257 6378
rect 4291 6344 4325 6378
rect 4359 6344 4393 6378
rect 4427 6344 4461 6378
rect 4495 6344 4529 6378
rect 4563 6344 4597 6378
rect 4631 6344 4665 6378
rect 4699 6344 4733 6378
rect 4767 6344 4801 6378
rect 4835 6344 4869 6378
rect 4903 6344 4937 6378
rect 4971 6344 5005 6378
rect 5039 6344 5073 6378
rect 5107 6349 5584 6378
rect 5904 6377 5945 6411
rect 5979 6377 6020 6411
rect 6054 6377 6095 6411
rect 6129 6377 6170 6411
rect 6204 6377 6245 6411
rect 6279 6377 6319 6411
rect 6353 6377 6393 6411
rect 5107 6344 5180 6349
rect 3340 6315 5180 6344
rect 5214 6315 5248 6349
rect 5282 6315 5316 6349
rect 5350 6315 5384 6349
rect 5418 6315 5452 6349
rect 5486 6315 5520 6349
rect 5554 6315 5584 6349
rect 3340 6308 5584 6315
rect 3340 6274 3373 6308
rect 3407 6274 3441 6308
rect 3475 6274 3509 6308
rect 3543 6274 3577 6308
rect 3611 6274 3645 6308
rect 3679 6274 3713 6308
rect 3747 6274 3781 6308
rect 3815 6274 3849 6308
rect 3883 6274 3917 6308
rect 3951 6274 3985 6308
rect 4019 6274 4053 6308
rect 4087 6274 4121 6308
rect 4155 6274 4189 6308
rect 4223 6274 4257 6308
rect 4291 6274 4325 6308
rect 4359 6274 4393 6308
rect 4427 6274 4461 6308
rect 4495 6274 4529 6308
rect 4563 6274 4597 6308
rect 4631 6274 4665 6308
rect 4699 6274 4733 6308
rect 4767 6274 4801 6308
rect 4835 6274 4869 6308
rect 4903 6274 4937 6308
rect 4971 6274 5005 6308
rect 5039 6274 5073 6308
rect 5107 6274 5584 6308
rect 3340 6242 5584 6274
rect 6852 6281 6886 6295
rect 6966 6289 7005 6323
rect 7039 6289 7078 6323
rect 7112 6289 7151 6323
rect 7185 6289 7224 6323
rect 7258 6289 7297 6323
rect 7331 6289 7370 6323
rect 7404 6289 7443 6323
rect 7477 6289 7516 6323
rect 7550 6289 7589 6323
rect 7623 6289 7662 6323
rect 7696 6289 7735 6323
rect 7769 6289 7808 6323
rect 7842 6289 7881 6323
rect 7915 6289 7954 6323
rect 7988 6289 8027 6323
rect 8061 6289 8100 6323
rect 8134 6289 8173 6323
rect 8207 6289 8246 6323
rect 8280 6289 8319 6323
rect 8353 6289 8392 6323
rect 8426 6289 8465 6323
rect 8499 6289 8538 6323
rect 8572 6289 8611 6323
rect 8645 6289 8684 6323
rect 8718 6289 8757 6323
rect 8791 6289 8830 6323
rect 8864 6289 8903 6323
rect 8937 6289 8976 6323
rect 9010 6289 9049 6323
rect 9083 6289 9122 6323
rect 9156 6289 9195 6323
rect 9229 6289 9268 6323
rect 9302 6289 9341 6323
rect 9375 6289 9414 6323
rect 9448 6289 9486 6323
rect 9520 6289 9558 6323
rect 9592 6289 9630 6323
rect 9664 6289 9702 6323
rect 9736 6289 9774 6323
rect 9808 6289 9846 6323
rect 10165 6289 10203 6323
rect 10237 6289 10275 6323
rect 10309 6289 10347 6323
rect 10381 6289 10419 6323
rect 10453 6289 10491 6323
rect 10525 6289 10563 6323
rect 10597 6289 10635 6323
rect 10669 6289 10707 6323
rect 10741 6289 10779 6323
rect 10813 6289 10852 6323
rect 10886 6289 10925 6323
rect 10959 6289 10998 6323
rect 11032 6289 11071 6323
rect 11105 6289 11144 6323
rect 11178 6289 11217 6323
rect 11251 6289 11290 6323
rect 11324 6289 11363 6323
rect 11397 6289 11436 6323
rect 11470 6289 11509 6323
rect 11543 6289 11582 6323
rect 11616 6289 11655 6323
rect 11689 6289 11728 6323
rect 11762 6289 11801 6323
rect 11835 6289 11874 6323
rect 11908 6289 11947 6323
rect 11981 6289 12020 6323
rect 12054 6289 12093 6323
rect 12127 6289 12166 6323
rect 12200 6289 12239 6323
rect 12273 6289 12312 6323
rect 12346 6289 12385 6323
rect 12419 6289 12458 6323
rect 12492 6289 12531 6323
rect 12565 6289 12604 6323
rect 12638 6289 12677 6323
rect 12711 6289 12750 6323
rect 12784 6289 12823 6323
rect 12857 6289 12896 6323
rect 12930 6289 12969 6323
rect 13003 6289 13042 6323
rect 13125 6281 13159 6295
rect 3340 6238 6781 6242
rect 3340 6204 3373 6238
rect 3407 6204 3441 6238
rect 3475 6204 3509 6238
rect 3543 6204 3577 6238
rect 3611 6204 3645 6238
rect 3679 6204 3713 6238
rect 3747 6204 3781 6238
rect 3815 6204 3849 6238
rect 3883 6204 3917 6238
rect 3951 6204 3985 6238
rect 4019 6204 4053 6238
rect 4087 6204 4121 6238
rect 4155 6204 4189 6238
rect 4223 6204 4257 6238
rect 4291 6204 4325 6238
rect 4359 6204 4393 6238
rect 4427 6204 4461 6238
rect 4495 6204 4529 6238
rect 4563 6204 4597 6238
rect 4631 6204 4665 6238
rect 4699 6204 4733 6238
rect 4767 6204 4801 6238
rect 4835 6204 4869 6238
rect 4903 6204 4937 6238
rect 4971 6204 5005 6238
rect 5039 6204 5073 6238
rect 5107 6218 6781 6238
rect 5107 6204 5155 6218
rect 3340 6184 5155 6204
rect 5189 6184 5223 6218
rect 5257 6184 5291 6218
rect 5325 6184 5359 6218
rect 5393 6184 5427 6218
rect 5461 6184 5495 6218
rect 5529 6184 5563 6218
rect 5597 6184 5631 6218
rect 5665 6184 5699 6218
rect 5733 6184 5767 6218
rect 5801 6184 5835 6218
rect 5869 6184 5903 6218
rect 5937 6184 5971 6218
rect 6005 6184 6040 6218
rect 6074 6184 6108 6218
rect 6142 6184 6176 6218
rect 6210 6184 6244 6218
rect 6278 6184 6312 6218
rect 6346 6184 6380 6218
rect 6414 6184 6448 6218
rect 6482 6184 6516 6218
rect 6550 6184 6584 6218
rect 6618 6184 6652 6218
rect 6686 6184 6720 6218
rect 6754 6184 6781 6218
rect 3340 6168 6781 6184
rect 3340 6134 3373 6168
rect 3407 6134 3441 6168
rect 3475 6134 3509 6168
rect 3543 6134 3577 6168
rect 3611 6134 3645 6168
rect 3679 6134 3713 6168
rect 3747 6134 3781 6168
rect 3815 6134 3849 6168
rect 3883 6134 3917 6168
rect 3951 6134 3985 6168
rect 4019 6134 4053 6168
rect 4087 6134 4121 6168
rect 4155 6134 4189 6168
rect 4223 6134 4257 6168
rect 4291 6134 4325 6168
rect 4359 6134 4393 6168
rect 4427 6134 4461 6168
rect 4495 6134 4529 6168
rect 4563 6134 4597 6168
rect 4631 6134 4665 6168
rect 4699 6134 4733 6168
rect 4767 6134 4801 6168
rect 4835 6134 4869 6168
rect 4903 6134 4937 6168
rect 4971 6134 5005 6168
rect 5039 6134 5073 6168
rect 5107 6149 6781 6168
rect 6852 6211 6886 6245
rect 13156 6279 13159 6281
rect 13122 6245 13125 6247
rect 13122 6211 13159 6245
rect 13122 6209 13125 6211
rect 13156 6175 13159 6177
rect 6852 6161 6886 6175
rect 5107 6148 6040 6149
rect 5107 6134 5155 6148
rect 3340 6114 5155 6134
rect 5189 6114 5223 6148
rect 5257 6114 5291 6148
rect 5325 6114 5359 6148
rect 5393 6114 5427 6148
rect 5461 6114 5495 6148
rect 5529 6114 5563 6148
rect 5597 6114 5631 6148
rect 5665 6114 5699 6148
rect 5733 6114 5767 6148
rect 5801 6114 5835 6148
rect 5869 6114 5903 6148
rect 5937 6114 5971 6148
rect 6005 6115 6040 6148
rect 6074 6115 6108 6149
rect 6142 6115 6176 6149
rect 6210 6115 6244 6149
rect 6278 6115 6312 6149
rect 6346 6115 6380 6149
rect 6414 6115 6448 6149
rect 6482 6115 6516 6149
rect 6550 6115 6584 6149
rect 6618 6115 6652 6149
rect 6686 6115 6720 6149
rect 6754 6115 6781 6149
rect 7206 6133 7246 6167
rect 7280 6133 7320 6167
rect 7354 6133 7394 6167
rect 7428 6133 7468 6167
rect 7502 6133 7542 6167
rect 7576 6133 7616 6167
rect 7650 6133 7690 6167
rect 7724 6133 7764 6167
rect 7798 6133 7837 6167
rect 7871 6133 7910 6167
rect 7944 6133 7983 6167
rect 8017 6133 8056 6167
rect 8090 6133 8129 6167
rect 8163 6133 8202 6167
rect 8236 6133 8275 6167
rect 8309 6133 8348 6167
rect 8382 6133 8421 6167
rect 8455 6133 8494 6167
rect 8528 6133 8567 6167
rect 8601 6133 8640 6167
rect 8674 6133 8713 6167
rect 8747 6133 8786 6167
rect 8820 6133 8859 6167
rect 8893 6133 8932 6167
rect 8966 6133 9005 6167
rect 9039 6133 9078 6167
rect 9112 6133 9151 6167
rect 9185 6133 9224 6167
rect 9258 6133 9297 6167
rect 9331 6133 9370 6167
rect 9404 6133 9443 6167
rect 9477 6133 9516 6167
rect 9550 6133 9589 6167
rect 9623 6133 9662 6167
rect 9696 6133 9735 6167
rect 9769 6133 9808 6167
rect 10203 6133 10242 6167
rect 10276 6133 10315 6167
rect 10349 6133 10388 6167
rect 10422 6133 10461 6167
rect 10495 6133 10534 6167
rect 10568 6133 10607 6167
rect 10641 6133 10680 6167
rect 10714 6133 10753 6167
rect 10787 6133 10826 6167
rect 10860 6133 10899 6167
rect 10933 6133 10972 6167
rect 11006 6133 11045 6167
rect 11079 6133 11118 6167
rect 11152 6133 11191 6167
rect 11225 6133 11264 6167
rect 11298 6133 11337 6167
rect 11371 6133 11410 6167
rect 11444 6133 11483 6167
rect 11517 6133 11556 6167
rect 11590 6133 11629 6167
rect 11663 6133 11702 6167
rect 11736 6133 11775 6167
rect 11809 6133 11848 6167
rect 11882 6133 11921 6167
rect 11955 6133 11994 6167
rect 12028 6133 12067 6167
rect 12101 6133 12140 6167
rect 12174 6133 12213 6167
rect 12247 6133 12286 6167
rect 12320 6133 12359 6167
rect 12393 6133 12432 6167
rect 12466 6133 12506 6167
rect 12540 6133 12580 6167
rect 12614 6133 12654 6167
rect 12688 6133 12728 6167
rect 12762 6133 12802 6167
rect 13125 6161 13159 6175
rect 6005 6114 6781 6115
rect 3340 6098 6781 6114
rect 3340 6064 3373 6098
rect 3407 6064 3441 6098
rect 3475 6064 3509 6098
rect 3543 6064 3577 6098
rect 3611 6064 3645 6098
rect 3679 6064 3713 6098
rect 3747 6064 3781 6098
rect 3815 6064 3849 6098
rect 3883 6064 3917 6098
rect 3951 6064 3985 6098
rect 4019 6064 4053 6098
rect 4087 6064 4121 6098
rect 4155 6064 4189 6098
rect 4223 6064 4257 6098
rect 4291 6064 4325 6098
rect 4359 6064 4393 6098
rect 4427 6064 4461 6098
rect 4495 6064 4529 6098
rect 4563 6064 4597 6098
rect 4631 6064 4665 6098
rect 4699 6064 4733 6098
rect 4767 6064 4801 6098
rect 4835 6064 4869 6098
rect 4903 6064 4937 6098
rect 4971 6064 5005 6098
rect 5039 6064 5073 6098
rect 5107 6080 6781 6098
rect 5107 6078 6040 6080
rect 5107 6064 5155 6078
rect 3340 6044 5155 6064
rect 5189 6044 5223 6078
rect 5257 6044 5291 6078
rect 5325 6044 5359 6078
rect 5393 6044 5427 6078
rect 5461 6044 5495 6078
rect 5529 6044 5563 6078
rect 5597 6044 5631 6078
rect 5665 6044 5699 6078
rect 5733 6044 5767 6078
rect 5801 6044 5835 6078
rect 5869 6044 5903 6078
rect 5937 6044 5971 6078
rect 6005 6046 6040 6078
rect 6074 6046 6108 6080
rect 6142 6046 6176 6080
rect 6210 6046 6244 6080
rect 6278 6046 6312 6080
rect 6346 6046 6380 6080
rect 6414 6046 6448 6080
rect 6482 6046 6516 6080
rect 6550 6046 6584 6080
rect 6618 6046 6652 6080
rect 6686 6046 6720 6080
rect 6754 6071 6781 6080
rect 6754 6046 6825 6071
rect 6005 6044 6825 6046
rect 3340 6037 6825 6044
rect 6859 6037 6893 6071
rect 6927 6037 6961 6071
rect 6995 6037 7029 6071
rect 7063 6037 7097 6071
rect 7131 6037 7165 6071
rect 7199 6037 7233 6071
rect 7267 6037 7301 6071
rect 7335 6037 7369 6071
rect 7403 6037 7437 6071
rect 7471 6037 7505 6071
rect 7539 6037 7573 6071
rect 7607 6037 7641 6071
rect 7675 6037 7709 6071
rect 7743 6037 7777 6071
rect 7811 6037 7845 6071
rect 7879 6037 7913 6071
rect 7947 6037 7981 6071
rect 8015 6037 8049 6071
rect 8083 6037 8117 6071
rect 8151 6037 8185 6071
rect 8219 6037 8253 6071
rect 8287 6037 8321 6071
rect 8355 6037 8389 6071
rect 8423 6037 8457 6071
rect 8491 6037 8525 6071
rect 8559 6037 8593 6071
rect 8627 6037 8661 6071
rect 8695 6037 8729 6071
rect 8763 6037 8797 6071
rect 8831 6037 8865 6071
rect 8899 6037 8933 6071
rect 8967 6037 9001 6071
rect 9035 6037 9069 6071
rect 9103 6037 9137 6071
rect 9171 6037 9205 6071
rect 9239 6037 9273 6071
rect 9307 6037 9341 6071
rect 9375 6037 9409 6071
rect 9443 6037 9477 6071
rect 9511 6037 9545 6071
rect 9579 6037 9613 6071
rect 9647 6037 9681 6071
rect 9715 6037 9749 6071
rect 9783 6037 9817 6071
rect 9851 6037 9886 6071
rect 9920 6037 9955 6071
rect 9989 6037 10024 6071
rect 10058 6037 10093 6071
rect 10127 6037 10162 6071
rect 10196 6037 10231 6071
rect 10265 6037 10300 6071
rect 10334 6037 10369 6071
rect 10403 6037 10438 6071
rect 10472 6037 10507 6071
rect 10541 6037 10576 6071
rect 10610 6037 10645 6071
rect 10679 6037 10714 6071
rect 10748 6037 10783 6071
rect 10817 6037 10852 6071
rect 10886 6037 10921 6071
rect 10955 6037 10990 6071
rect 11024 6037 11059 6071
rect 11093 6037 11128 6071
rect 11162 6037 11197 6071
rect 11231 6037 11266 6071
rect 11300 6037 11335 6071
rect 11369 6037 11404 6071
rect 11438 6037 11473 6071
rect 11507 6037 11542 6071
rect 11576 6037 11611 6071
rect 11645 6037 11680 6071
rect 11714 6037 11749 6071
rect 11783 6037 11818 6071
rect 11852 6037 11887 6071
rect 11921 6037 11956 6071
rect 11990 6037 12025 6071
rect 12059 6037 12094 6071
rect 12128 6037 12163 6071
rect 12197 6037 12232 6071
rect 12266 6037 12301 6071
rect 12335 6037 12370 6071
rect 12404 6037 12439 6071
rect 12473 6037 12508 6071
rect 12542 6037 12577 6071
rect 12611 6037 12646 6071
rect 12680 6037 12715 6071
rect 12749 6037 12784 6071
rect 12818 6037 12853 6071
rect 12887 6037 12922 6071
rect 12956 6037 12991 6071
rect 13025 6037 13060 6071
rect 13094 6037 13129 6071
rect 13163 6037 13197 6071
rect 3340 6028 6781 6037
rect 3340 5994 3373 6028
rect 3407 5994 3441 6028
rect 3475 5994 3509 6028
rect 3543 5994 3577 6028
rect 3611 5994 3645 6028
rect 3679 5994 3713 6028
rect 3747 5994 3781 6028
rect 3815 5994 3849 6028
rect 3883 5994 3917 6028
rect 3951 5994 3985 6028
rect 4019 5994 4053 6028
rect 4087 5994 4121 6028
rect 4155 5994 4189 6028
rect 4223 5994 4257 6028
rect 4291 5994 4325 6028
rect 4359 5994 4393 6028
rect 4427 5994 4461 6028
rect 4495 5994 4529 6028
rect 4563 5994 4597 6028
rect 4631 5994 4665 6028
rect 4699 5994 4733 6028
rect 4767 5994 4801 6028
rect 4835 5994 4869 6028
rect 4903 5994 4937 6028
rect 4971 5994 5005 6028
rect 5039 5994 5073 6028
rect 5107 6011 6781 6028
rect 5107 6008 6040 6011
rect 5107 5994 5155 6008
rect 3340 5974 5155 5994
rect 5189 5974 5223 6008
rect 5257 5974 5291 6008
rect 5325 5974 5359 6008
rect 5393 5974 5427 6008
rect 5461 5974 5495 6008
rect 5529 5974 5563 6008
rect 5597 5974 5631 6008
rect 5665 5974 5699 6008
rect 5733 5974 5767 6008
rect 5801 5974 5835 6008
rect 5869 5974 5903 6008
rect 5937 5974 5971 6008
rect 6005 5977 6040 6008
rect 6074 5977 6108 6011
rect 6142 5977 6176 6011
rect 6210 5977 6244 6011
rect 6278 5977 6312 6011
rect 6346 5977 6380 6011
rect 6414 5977 6448 6011
rect 6482 5977 6516 6011
rect 6550 5977 6584 6011
rect 6618 5977 6652 6011
rect 6686 5977 6720 6011
rect 6754 5977 6781 6011
rect 6005 5974 6781 5977
rect 3340 5958 6781 5974
rect 3340 5924 3373 5958
rect 3407 5924 3441 5958
rect 3475 5924 3509 5958
rect 3543 5924 3577 5958
rect 3611 5924 3645 5958
rect 3679 5924 3713 5958
rect 3747 5924 3781 5958
rect 3815 5924 3849 5958
rect 3883 5924 3917 5958
rect 3951 5924 3985 5958
rect 4019 5924 4053 5958
rect 4087 5924 4121 5958
rect 4155 5924 4189 5958
rect 4223 5924 4257 5958
rect 4291 5924 4325 5958
rect 4359 5924 4393 5958
rect 4427 5924 4461 5958
rect 4495 5924 4529 5958
rect 4563 5924 4597 5958
rect 4631 5924 4665 5958
rect 4699 5924 4733 5958
rect 4767 5924 4801 5958
rect 4835 5924 4869 5958
rect 4903 5924 4937 5958
rect 4971 5924 5005 5958
rect 5039 5924 5073 5958
rect 5107 5942 6781 5958
rect 5107 5938 6040 5942
rect 5107 5924 5155 5938
rect 3340 5904 5155 5924
rect 5189 5904 5223 5938
rect 5257 5904 5291 5938
rect 5325 5904 5359 5938
rect 5393 5904 5427 5938
rect 5461 5904 5495 5938
rect 5529 5904 5563 5938
rect 5597 5904 5631 5938
rect 5665 5904 5699 5938
rect 5733 5904 5767 5938
rect 5801 5904 5835 5938
rect 5869 5904 5903 5938
rect 5937 5904 5971 5938
rect 6005 5908 6040 5938
rect 6074 5908 6108 5942
rect 6142 5908 6176 5942
rect 6210 5908 6244 5942
rect 6278 5908 6312 5942
rect 6346 5908 6380 5942
rect 6414 5908 6448 5942
rect 6482 5908 6516 5942
rect 6550 5908 6584 5942
rect 6618 5908 6652 5942
rect 6686 5908 6720 5942
rect 6754 5908 6781 5942
rect 6005 5904 6781 5908
rect 3340 5888 6781 5904
rect 3340 5854 3373 5888
rect 3407 5854 3441 5888
rect 3475 5854 3509 5888
rect 3543 5854 3577 5888
rect 3611 5854 3645 5888
rect 3679 5854 3713 5888
rect 3747 5854 3781 5888
rect 3815 5854 3849 5888
rect 3883 5854 3917 5888
rect 3951 5854 3985 5888
rect 4019 5854 4053 5888
rect 4087 5854 4121 5888
rect 4155 5854 4189 5888
rect 4223 5854 4257 5888
rect 4291 5854 4325 5888
rect 4359 5854 4393 5888
rect 4427 5854 4461 5888
rect 4495 5854 4529 5888
rect 4563 5854 4597 5888
rect 4631 5854 4665 5888
rect 4699 5854 4733 5888
rect 4767 5854 4801 5888
rect 4835 5854 4869 5888
rect 4903 5854 4937 5888
rect 4971 5854 5005 5888
rect 5039 5854 5073 5888
rect 5107 5873 6781 5888
rect 5107 5868 6040 5873
rect 5107 5854 5155 5868
rect 3340 5834 5155 5854
rect 5189 5834 5223 5868
rect 5257 5834 5291 5868
rect 5325 5834 5359 5868
rect 5393 5834 5427 5868
rect 5461 5834 5495 5868
rect 5529 5834 5563 5868
rect 5597 5834 5631 5868
rect 5665 5834 5699 5868
rect 5733 5834 5767 5868
rect 5801 5834 5835 5868
rect 5869 5834 5903 5868
rect 5937 5834 5971 5868
rect 6005 5839 6040 5868
rect 6074 5839 6108 5873
rect 6142 5839 6176 5873
rect 6210 5839 6244 5873
rect 6278 5839 6312 5873
rect 6346 5839 6380 5873
rect 6414 5839 6448 5873
rect 6482 5839 6516 5873
rect 6550 5839 6584 5873
rect 6618 5839 6652 5873
rect 6686 5839 6720 5873
rect 6754 5839 6781 5873
rect 6005 5834 6781 5839
rect 3340 5818 6781 5834
rect 3340 5784 3373 5818
rect 3407 5784 3441 5818
rect 3475 5784 3509 5818
rect 3543 5784 3577 5818
rect 3611 5784 3645 5818
rect 3679 5784 3713 5818
rect 3747 5784 3781 5818
rect 3815 5784 3849 5818
rect 3883 5784 3917 5818
rect 3951 5784 3985 5818
rect 4019 5784 4053 5818
rect 4087 5784 4121 5818
rect 4155 5784 4189 5818
rect 4223 5784 4257 5818
rect 4291 5784 4325 5818
rect 4359 5784 4393 5818
rect 4427 5784 4461 5818
rect 4495 5784 4529 5818
rect 4563 5784 4597 5818
rect 4631 5784 4665 5818
rect 4699 5784 4733 5818
rect 4767 5784 4801 5818
rect 4835 5784 4869 5818
rect 4903 5784 4937 5818
rect 4971 5784 5005 5818
rect 5039 5784 5073 5818
rect 5107 5804 6781 5818
rect 6852 5931 6886 5946
rect 6966 5941 7005 5975
rect 7039 5941 7078 5975
rect 7112 5941 7151 5975
rect 7185 5941 7224 5975
rect 7258 5941 7297 5975
rect 7331 5941 7370 5975
rect 7404 5941 7443 5975
rect 7477 5941 7516 5975
rect 7550 5941 7589 5975
rect 7623 5941 7662 5975
rect 7696 5941 7735 5975
rect 7769 5941 7808 5975
rect 7842 5941 7881 5975
rect 7915 5941 7954 5975
rect 7988 5941 8027 5975
rect 8061 5941 8100 5975
rect 8134 5941 8173 5975
rect 8207 5941 8246 5975
rect 8280 5941 8319 5975
rect 8353 5941 8392 5975
rect 8426 5941 8465 5975
rect 8499 5941 8538 5975
rect 8572 5941 8611 5975
rect 8645 5941 8684 5975
rect 8718 5941 8757 5975
rect 8791 5941 8830 5975
rect 8864 5941 8903 5975
rect 8937 5941 8976 5975
rect 9010 5941 9049 5975
rect 9083 5941 9122 5975
rect 9156 5941 9195 5975
rect 9229 5941 9268 5975
rect 9302 5941 9341 5975
rect 9375 5941 9414 5975
rect 9448 5941 9486 5975
rect 9520 5941 9558 5975
rect 9592 5941 9630 5975
rect 9664 5941 9702 5975
rect 9736 5941 9774 5975
rect 9808 5941 9846 5975
rect 10165 5941 10203 5975
rect 10237 5941 10275 5975
rect 10309 5941 10347 5975
rect 10381 5941 10419 5975
rect 10453 5941 10491 5975
rect 10525 5941 10563 5975
rect 10597 5941 10635 5975
rect 10669 5941 10707 5975
rect 10741 5941 10779 5975
rect 10813 5941 10852 5975
rect 10886 5941 10925 5975
rect 10959 5941 10998 5975
rect 11032 5941 11071 5975
rect 11105 5941 11144 5975
rect 11178 5941 11217 5975
rect 11251 5941 11290 5975
rect 11324 5941 11363 5975
rect 11397 5941 11436 5975
rect 11470 5941 11509 5975
rect 11543 5941 11582 5975
rect 11616 5941 11655 5975
rect 11689 5941 11728 5975
rect 11762 5941 11801 5975
rect 11835 5941 11874 5975
rect 11908 5941 11947 5975
rect 11981 5941 12020 5975
rect 12054 5941 12093 5975
rect 12127 5941 12166 5975
rect 12200 5941 12239 5975
rect 12273 5941 12312 5975
rect 12346 5941 12385 5975
rect 12419 5941 12458 5975
rect 12492 5941 12531 5975
rect 12565 5941 12604 5975
rect 12638 5941 12677 5975
rect 12711 5941 12750 5975
rect 12784 5941 12823 5975
rect 12857 5941 12896 5975
rect 12930 5941 12969 5975
rect 13003 5941 13042 5975
rect 13125 5933 13159 5947
rect 6852 5862 6886 5896
rect 13156 5931 13159 5933
rect 13122 5897 13125 5899
rect 13122 5863 13159 5897
rect 13122 5861 13125 5863
rect 13156 5827 13159 5829
rect 6852 5812 6886 5825
rect 5107 5798 6040 5804
rect 5107 5784 5155 5798
rect 3340 5764 5155 5784
rect 5189 5764 5223 5798
rect 5257 5764 5291 5798
rect 5325 5764 5359 5798
rect 5393 5764 5427 5798
rect 5461 5764 5495 5798
rect 5529 5764 5563 5798
rect 5597 5764 5631 5798
rect 5665 5764 5699 5798
rect 5733 5764 5767 5798
rect 5801 5764 5835 5798
rect 5869 5764 5903 5798
rect 5937 5764 5971 5798
rect 6005 5770 6040 5798
rect 6074 5770 6108 5804
rect 6142 5770 6176 5804
rect 6210 5770 6244 5804
rect 6278 5770 6312 5804
rect 6346 5770 6380 5804
rect 6414 5770 6448 5804
rect 6482 5770 6516 5804
rect 6550 5770 6584 5804
rect 6618 5770 6652 5804
rect 6686 5770 6720 5804
rect 6754 5770 6781 5804
rect 7215 5785 7254 5819
rect 7288 5785 7327 5819
rect 7361 5785 7400 5819
rect 7434 5785 7473 5819
rect 7507 5785 7546 5819
rect 7580 5785 7619 5819
rect 7653 5785 7692 5819
rect 7726 5785 7765 5819
rect 7799 5785 7838 5819
rect 7872 5785 7911 5819
rect 7945 5785 7984 5819
rect 8018 5785 8057 5819
rect 8091 5785 8130 5819
rect 8164 5785 8203 5819
rect 8237 5785 8276 5819
rect 8310 5785 8349 5819
rect 8383 5785 8422 5819
rect 8456 5785 8494 5819
rect 8528 5785 8566 5819
rect 8600 5785 8638 5819
rect 8672 5785 8710 5819
rect 8744 5785 8782 5819
rect 8816 5785 8854 5819
rect 8888 5785 8926 5819
rect 8960 5785 8998 5819
rect 9032 5785 9070 5819
rect 9104 5785 9142 5819
rect 9176 5785 9214 5819
rect 9248 5785 9286 5819
rect 9320 5785 9358 5819
rect 9392 5785 9430 5819
rect 9464 5785 9502 5819
rect 9536 5785 9574 5819
rect 10203 5785 10242 5819
rect 10276 5785 10315 5819
rect 10349 5785 10388 5819
rect 10422 5785 10461 5819
rect 10495 5785 10534 5819
rect 10568 5785 10607 5819
rect 10641 5785 10680 5819
rect 10714 5785 10753 5819
rect 10787 5785 10826 5819
rect 10860 5785 10899 5819
rect 10933 5785 10972 5819
rect 11006 5785 11045 5819
rect 11079 5785 11118 5819
rect 11152 5785 11191 5819
rect 11225 5785 11264 5819
rect 11298 5785 11337 5819
rect 11371 5785 11410 5819
rect 11444 5785 11483 5819
rect 11517 5785 11556 5819
rect 11590 5785 11629 5819
rect 11663 5785 11702 5819
rect 11736 5785 11775 5819
rect 11809 5785 11848 5819
rect 11882 5785 11921 5819
rect 11955 5785 11994 5819
rect 12028 5785 12067 5819
rect 12101 5785 12140 5819
rect 12174 5785 12213 5819
rect 12247 5785 12286 5819
rect 12320 5785 12359 5819
rect 12393 5785 12432 5819
rect 12466 5785 12506 5819
rect 12540 5785 12580 5819
rect 12614 5785 12654 5819
rect 12688 5785 12728 5819
rect 12762 5785 12802 5819
rect 13125 5813 13159 5827
rect 6005 5764 6781 5770
rect 3340 5748 6781 5764
rect 3340 5714 3373 5748
rect 3407 5714 3441 5748
rect 3475 5714 3509 5748
rect 3543 5714 3577 5748
rect 3611 5714 3645 5748
rect 3679 5714 3713 5748
rect 3747 5714 3781 5748
rect 3815 5714 3849 5748
rect 3883 5714 3917 5748
rect 3951 5714 3985 5748
rect 4019 5714 4053 5748
rect 4087 5714 4121 5748
rect 4155 5714 4189 5748
rect 4223 5714 4257 5748
rect 4291 5714 4325 5748
rect 4359 5714 4393 5748
rect 4427 5714 4461 5748
rect 4495 5714 4529 5748
rect 4563 5714 4597 5748
rect 4631 5714 4665 5748
rect 4699 5714 4733 5748
rect 4767 5714 4801 5748
rect 4835 5714 4869 5748
rect 4903 5714 4937 5748
rect 4971 5714 5005 5748
rect 5039 5714 5073 5748
rect 5107 5735 6781 5748
rect 5107 5728 6040 5735
rect 5107 5714 5155 5728
rect 3340 5694 5155 5714
rect 5189 5694 5223 5728
rect 5257 5694 5291 5728
rect 5325 5694 5359 5728
rect 5393 5694 5427 5728
rect 5461 5694 5495 5728
rect 5529 5694 5563 5728
rect 5597 5694 5631 5728
rect 5665 5694 5699 5728
rect 5733 5694 5767 5728
rect 5801 5694 5835 5728
rect 5869 5694 5903 5728
rect 5937 5694 5971 5728
rect 6005 5701 6040 5728
rect 6074 5701 6108 5735
rect 6142 5701 6176 5735
rect 6210 5701 6244 5735
rect 6278 5701 6312 5735
rect 6346 5701 6380 5735
rect 6414 5701 6448 5735
rect 6482 5701 6516 5735
rect 6550 5701 6584 5735
rect 6618 5701 6652 5735
rect 6686 5701 6720 5735
rect 6754 5723 6781 5735
rect 6754 5701 6825 5723
rect 6005 5694 6825 5701
rect 3340 5689 6825 5694
rect 6859 5689 6893 5723
rect 6927 5689 6961 5723
rect 6995 5689 7029 5723
rect 7063 5689 7097 5723
rect 7131 5689 7165 5723
rect 7199 5689 7233 5723
rect 7267 5689 7301 5723
rect 7335 5689 7369 5723
rect 7403 5689 7437 5723
rect 7471 5689 7505 5723
rect 7539 5689 7573 5723
rect 7607 5689 7641 5723
rect 7675 5689 7709 5723
rect 7743 5689 7777 5723
rect 7811 5689 7845 5723
rect 7879 5689 7913 5723
rect 7947 5689 7981 5723
rect 8015 5689 8049 5723
rect 8083 5689 8117 5723
rect 8151 5689 8185 5723
rect 8219 5689 8253 5723
rect 8287 5689 8321 5723
rect 8355 5689 8389 5723
rect 8423 5689 8457 5723
rect 8491 5689 8525 5723
rect 8559 5689 8593 5723
rect 8627 5689 8661 5723
rect 8695 5689 8729 5723
rect 8763 5689 8797 5723
rect 8831 5689 8865 5723
rect 8899 5689 8933 5723
rect 8967 5689 9001 5723
rect 9035 5689 9069 5723
rect 9103 5689 9137 5723
rect 9171 5689 9205 5723
rect 9239 5689 9273 5723
rect 9307 5689 9341 5723
rect 9375 5689 9409 5723
rect 9443 5689 9477 5723
rect 9511 5689 9545 5723
rect 9579 5689 9613 5723
rect 9647 5689 9681 5723
rect 9715 5689 9749 5723
rect 9783 5689 9817 5723
rect 9851 5689 9886 5723
rect 9920 5689 9955 5723
rect 9989 5689 10024 5723
rect 10058 5689 10093 5723
rect 10127 5689 10162 5723
rect 10196 5689 10231 5723
rect 10265 5689 10300 5723
rect 10334 5689 10369 5723
rect 10403 5689 10438 5723
rect 10472 5689 10507 5723
rect 10541 5689 10576 5723
rect 10610 5689 10645 5723
rect 10679 5689 10714 5723
rect 10748 5689 10783 5723
rect 10817 5689 10852 5723
rect 10886 5689 10921 5723
rect 10955 5689 10990 5723
rect 11024 5689 11059 5723
rect 11093 5689 11128 5723
rect 11162 5689 11197 5723
rect 11231 5689 11266 5723
rect 11300 5689 11335 5723
rect 11369 5689 11404 5723
rect 11438 5689 11473 5723
rect 11507 5689 11542 5723
rect 11576 5689 11611 5723
rect 11645 5689 11680 5723
rect 11714 5689 11749 5723
rect 11783 5689 11818 5723
rect 11852 5689 11887 5723
rect 11921 5689 11956 5723
rect 11990 5689 12025 5723
rect 12059 5689 12094 5723
rect 12128 5689 12163 5723
rect 12197 5689 12232 5723
rect 12266 5689 12301 5723
rect 12335 5689 12370 5723
rect 12404 5689 12439 5723
rect 12473 5689 12508 5723
rect 12542 5689 12577 5723
rect 12611 5689 12646 5723
rect 12680 5689 12715 5723
rect 12749 5689 12784 5723
rect 12818 5689 12853 5723
rect 12887 5689 12922 5723
rect 12956 5689 12991 5723
rect 13025 5689 13060 5723
rect 13094 5689 13129 5723
rect 13163 5689 13197 5723
rect 3340 5678 6781 5689
rect 3340 5644 3373 5678
rect 3407 5644 3441 5678
rect 3475 5644 3509 5678
rect 3543 5644 3577 5678
rect 3611 5644 3645 5678
rect 3679 5644 3713 5678
rect 3747 5644 3781 5678
rect 3815 5644 3849 5678
rect 3883 5644 3917 5678
rect 3951 5644 3985 5678
rect 4019 5644 4053 5678
rect 4087 5644 4121 5678
rect 4155 5644 4189 5678
rect 4223 5644 4257 5678
rect 4291 5644 4325 5678
rect 4359 5644 4393 5678
rect 4427 5644 4461 5678
rect 4495 5644 4529 5678
rect 4563 5644 4597 5678
rect 4631 5644 4665 5678
rect 4699 5644 4733 5678
rect 4767 5644 4801 5678
rect 4835 5644 4869 5678
rect 4903 5644 4937 5678
rect 4971 5644 5005 5678
rect 5039 5644 5073 5678
rect 5107 5666 6781 5678
rect 5107 5657 6040 5666
rect 5107 5644 5155 5657
rect 3340 5623 5155 5644
rect 5189 5623 5223 5657
rect 5257 5623 5291 5657
rect 5325 5623 5359 5657
rect 5393 5623 5427 5657
rect 5461 5623 5495 5657
rect 5529 5623 5563 5657
rect 5597 5623 5631 5657
rect 5665 5623 5699 5657
rect 5733 5623 5767 5657
rect 5801 5623 5835 5657
rect 5869 5623 5903 5657
rect 5937 5623 5971 5657
rect 6005 5632 6040 5657
rect 6074 5632 6108 5666
rect 6142 5632 6176 5666
rect 6210 5632 6244 5666
rect 6278 5632 6312 5666
rect 6346 5632 6380 5666
rect 6414 5632 6448 5666
rect 6482 5632 6516 5666
rect 6550 5632 6584 5666
rect 6618 5632 6652 5666
rect 6686 5632 6720 5666
rect 6754 5632 6781 5666
rect 6005 5623 6781 5632
rect 3340 5608 6781 5623
rect 3340 5574 3373 5608
rect 3407 5574 3441 5608
rect 3475 5574 3509 5608
rect 3543 5574 3577 5608
rect 3611 5574 3645 5608
rect 3679 5574 3713 5608
rect 3747 5574 3781 5608
rect 3815 5574 3849 5608
rect 3883 5574 3917 5608
rect 3951 5574 3985 5608
rect 4019 5574 4053 5608
rect 4087 5574 4121 5608
rect 4155 5574 4189 5608
rect 4223 5574 4257 5608
rect 4291 5574 4325 5608
rect 4359 5574 4393 5608
rect 4427 5574 4461 5608
rect 4495 5574 4529 5608
rect 4563 5574 4597 5608
rect 4631 5574 4665 5608
rect 4699 5574 4733 5608
rect 4767 5574 4801 5608
rect 4835 5574 4869 5608
rect 4903 5574 4937 5608
rect 4971 5574 5005 5608
rect 5039 5574 5073 5608
rect 5107 5597 6781 5608
rect 5107 5586 6040 5597
rect 5107 5574 5155 5586
rect 3340 5552 5155 5574
rect 5189 5552 5223 5586
rect 5257 5552 5291 5586
rect 5325 5552 5359 5586
rect 5393 5552 5427 5586
rect 5461 5552 5495 5586
rect 5529 5552 5563 5586
rect 5597 5552 5631 5586
rect 5665 5552 5699 5586
rect 5733 5552 5767 5586
rect 5801 5552 5835 5586
rect 5869 5552 5903 5586
rect 5937 5552 5971 5586
rect 6005 5563 6040 5586
rect 6074 5563 6108 5597
rect 6142 5563 6176 5597
rect 6210 5563 6244 5597
rect 6278 5563 6312 5597
rect 6346 5563 6380 5597
rect 6414 5563 6448 5597
rect 6482 5563 6516 5597
rect 6550 5563 6584 5597
rect 6618 5563 6652 5597
rect 6686 5563 6720 5597
rect 6754 5563 6781 5597
rect 6005 5552 6781 5563
rect 3340 5538 6781 5552
rect 3340 5504 3373 5538
rect 3407 5504 3441 5538
rect 3475 5504 3509 5538
rect 3543 5504 3577 5538
rect 3611 5504 3645 5538
rect 3679 5504 3713 5538
rect 3747 5504 3781 5538
rect 3815 5504 3849 5538
rect 3883 5504 3917 5538
rect 3951 5504 3985 5538
rect 4019 5504 4053 5538
rect 4087 5504 4121 5538
rect 4155 5504 4189 5538
rect 4223 5504 4257 5538
rect 4291 5504 4325 5538
rect 4359 5504 4393 5538
rect 4427 5504 4461 5538
rect 4495 5504 4529 5538
rect 4563 5504 4597 5538
rect 4631 5504 4665 5538
rect 4699 5504 4733 5538
rect 4767 5504 4801 5538
rect 4835 5504 4869 5538
rect 4903 5504 4937 5538
rect 4971 5504 5005 5538
rect 5039 5504 5073 5538
rect 5107 5528 6781 5538
rect 5107 5505 6040 5528
rect 5107 5504 5155 5505
rect 3340 5471 5155 5504
rect 5189 5471 5223 5505
rect 5257 5471 5291 5505
rect 5325 5471 5359 5505
rect 5393 5471 5427 5505
rect 5461 5471 5495 5505
rect 5529 5471 5563 5505
rect 5597 5471 5631 5505
rect 5665 5471 5699 5505
rect 5733 5471 5767 5505
rect 5801 5471 5835 5505
rect 5869 5471 5903 5505
rect 5937 5471 5971 5505
rect 6005 5494 6040 5505
rect 6074 5494 6108 5528
rect 6142 5494 6176 5528
rect 6210 5494 6244 5528
rect 6278 5494 6312 5528
rect 6346 5494 6380 5528
rect 6414 5494 6448 5528
rect 6482 5494 6516 5528
rect 6550 5494 6584 5528
rect 6618 5494 6652 5528
rect 6686 5494 6720 5528
rect 6754 5494 6781 5528
rect 6005 5471 6781 5494
rect 3340 5468 6781 5471
rect 3340 5434 3373 5468
rect 3407 5434 3441 5468
rect 3475 5434 3509 5468
rect 3543 5434 3577 5468
rect 3611 5434 3645 5468
rect 3679 5434 3713 5468
rect 3747 5434 3781 5468
rect 3815 5434 3849 5468
rect 3883 5434 3917 5468
rect 3951 5434 3985 5468
rect 4019 5434 4053 5468
rect 4087 5434 4121 5468
rect 4155 5434 4189 5468
rect 4223 5434 4257 5468
rect 4291 5434 4325 5468
rect 4359 5434 4393 5468
rect 4427 5434 4461 5468
rect 4495 5434 4529 5468
rect 4563 5434 4597 5468
rect 4631 5434 4665 5468
rect 4699 5434 4733 5468
rect 4767 5434 4801 5468
rect 4835 5434 4869 5468
rect 4903 5434 4937 5468
rect 4971 5434 5005 5468
rect 5039 5434 5073 5468
rect 5107 5459 6781 5468
rect 6852 5584 6886 5599
rect 6966 5593 7005 5627
rect 7039 5593 7078 5627
rect 7112 5593 7151 5627
rect 7185 5593 7224 5627
rect 7258 5593 7297 5627
rect 7331 5593 7370 5627
rect 7404 5593 7443 5627
rect 7477 5593 7516 5627
rect 7550 5593 7589 5627
rect 7623 5593 7662 5627
rect 7696 5593 7735 5627
rect 7769 5593 7808 5627
rect 7842 5593 7881 5627
rect 7915 5593 7954 5627
rect 7988 5593 8027 5627
rect 8061 5593 8100 5627
rect 8134 5593 8173 5627
rect 8207 5593 8246 5627
rect 8280 5593 8319 5627
rect 8353 5593 8392 5627
rect 8426 5593 8465 5627
rect 8499 5593 8538 5627
rect 8572 5593 8611 5627
rect 8645 5593 8684 5627
rect 8718 5593 8757 5627
rect 8791 5593 8830 5627
rect 8864 5593 8903 5627
rect 8937 5593 8976 5627
rect 9010 5593 9049 5627
rect 9083 5593 9122 5627
rect 9156 5593 9195 5627
rect 9229 5593 9268 5627
rect 9302 5593 9341 5627
rect 9375 5593 9414 5627
rect 9448 5593 9486 5627
rect 9520 5593 9558 5627
rect 9592 5593 9630 5627
rect 9664 5593 9702 5627
rect 9736 5593 9774 5627
rect 9808 5593 9846 5627
rect 10165 5593 10203 5627
rect 10237 5593 10275 5627
rect 10309 5593 10347 5627
rect 10381 5593 10419 5627
rect 10453 5593 10491 5627
rect 10525 5593 10563 5627
rect 10597 5593 10635 5627
rect 10669 5593 10707 5627
rect 10741 5593 10779 5627
rect 10813 5593 10852 5627
rect 10886 5593 10925 5627
rect 10959 5593 10998 5627
rect 11032 5593 11071 5627
rect 11105 5593 11144 5627
rect 11178 5593 11217 5627
rect 11251 5593 11290 5627
rect 11324 5593 11363 5627
rect 11397 5593 11436 5627
rect 11470 5593 11509 5627
rect 11543 5593 11582 5627
rect 11616 5593 11655 5627
rect 11689 5593 11728 5627
rect 11762 5593 11801 5627
rect 11835 5593 11874 5627
rect 11908 5593 11947 5627
rect 11981 5593 12020 5627
rect 12054 5593 12093 5627
rect 12127 5593 12166 5627
rect 12200 5593 12239 5627
rect 12273 5593 12312 5627
rect 12346 5593 12385 5627
rect 12419 5593 12458 5627
rect 12492 5593 12531 5627
rect 12565 5593 12604 5627
rect 12638 5593 12677 5627
rect 12711 5593 12750 5627
rect 12784 5593 12823 5627
rect 12857 5593 12896 5627
rect 12930 5593 12969 5627
rect 13003 5593 13042 5627
rect 13125 5585 13159 5599
rect 6852 5515 6886 5549
rect 13156 5583 13159 5585
rect 13122 5549 13125 5551
rect 13122 5515 13159 5549
rect 13122 5513 13125 5515
rect 13156 5479 13159 5481
rect 6852 5465 6886 5478
rect 5107 5434 6040 5459
rect 3340 5431 6040 5434
rect 3340 5398 5155 5431
rect 3340 5364 3373 5398
rect 3407 5364 3441 5398
rect 3475 5364 3509 5398
rect 3543 5364 3577 5398
rect 3611 5364 3645 5398
rect 3679 5364 3713 5398
rect 3747 5364 3781 5398
rect 3815 5364 3849 5398
rect 3883 5364 3917 5398
rect 3951 5364 3985 5398
rect 4019 5364 4053 5398
rect 4087 5364 4121 5398
rect 4155 5364 4189 5398
rect 4223 5364 4257 5398
rect 4291 5364 4325 5398
rect 4359 5364 4393 5398
rect 4427 5364 4461 5398
rect 4495 5364 4529 5398
rect 4563 5364 4597 5398
rect 4631 5364 4665 5398
rect 4699 5364 4733 5398
rect 4767 5364 4801 5398
rect 4835 5364 4869 5398
rect 4903 5364 4937 5398
rect 4971 5364 5005 5398
rect 5039 5364 5073 5398
rect 5107 5397 5155 5398
rect 5189 5397 5223 5431
rect 5257 5397 5291 5431
rect 5325 5397 5359 5431
rect 5393 5397 5427 5431
rect 5461 5397 5495 5431
rect 5529 5397 5563 5431
rect 5597 5397 5631 5431
rect 5665 5397 5699 5431
rect 5733 5397 5767 5431
rect 5801 5397 5835 5431
rect 5869 5397 5903 5431
rect 5937 5397 5971 5431
rect 6005 5425 6040 5431
rect 6074 5425 6108 5459
rect 6142 5425 6176 5459
rect 6210 5425 6244 5459
rect 6278 5425 6312 5459
rect 6346 5425 6380 5459
rect 6414 5425 6448 5459
rect 6482 5425 6516 5459
rect 6550 5425 6584 5459
rect 6618 5425 6652 5459
rect 6686 5425 6720 5459
rect 6754 5425 6781 5459
rect 7206 5437 7246 5471
rect 7280 5437 7320 5471
rect 7354 5437 7394 5471
rect 7428 5437 7468 5471
rect 7502 5437 7542 5471
rect 7576 5437 7616 5471
rect 7650 5437 7690 5471
rect 7724 5437 7764 5471
rect 7798 5437 7838 5471
rect 7872 5437 7912 5471
rect 7946 5437 7985 5471
rect 8019 5437 8058 5471
rect 8092 5437 8131 5471
rect 8165 5437 8204 5471
rect 8238 5437 8277 5471
rect 8311 5437 8350 5471
rect 8384 5437 8423 5471
rect 8457 5437 8496 5471
rect 8530 5437 8569 5471
rect 8603 5437 8642 5471
rect 8676 5437 8715 5471
rect 8749 5437 8788 5471
rect 8822 5437 8861 5471
rect 8895 5437 8934 5471
rect 8968 5437 9007 5471
rect 9041 5437 9080 5471
rect 9114 5437 9153 5471
rect 9187 5437 9226 5471
rect 9260 5437 9299 5471
rect 9333 5437 9372 5471
rect 9406 5437 9445 5471
rect 9479 5437 9518 5471
rect 9552 5437 9591 5471
rect 9625 5437 9664 5471
rect 9698 5437 9737 5471
rect 9771 5437 9810 5471
rect 10203 5437 10242 5471
rect 10276 5437 10315 5471
rect 10349 5437 10388 5471
rect 10422 5437 10461 5471
rect 10495 5437 10534 5471
rect 10568 5437 10607 5471
rect 10641 5437 10680 5471
rect 10714 5437 10753 5471
rect 10787 5437 10826 5471
rect 10860 5437 10899 5471
rect 10933 5437 10972 5471
rect 11006 5437 11045 5471
rect 11079 5437 11118 5471
rect 11152 5437 11191 5471
rect 11225 5437 11264 5471
rect 11298 5437 11337 5471
rect 11371 5437 11410 5471
rect 11444 5437 11483 5471
rect 11517 5437 11556 5471
rect 11590 5437 11629 5471
rect 11663 5437 11702 5471
rect 11736 5437 11775 5471
rect 11809 5437 11848 5471
rect 11882 5437 11921 5471
rect 11955 5437 11994 5471
rect 12028 5437 12067 5471
rect 12101 5437 12140 5471
rect 12174 5437 12213 5471
rect 12247 5437 12286 5471
rect 12320 5437 12359 5471
rect 12393 5437 12432 5471
rect 12466 5437 12506 5471
rect 12540 5437 12580 5471
rect 12614 5437 12654 5471
rect 12688 5437 12728 5471
rect 12762 5437 12802 5471
rect 13125 5465 13159 5479
rect 6005 5397 6781 5425
rect 5107 5390 6781 5397
rect 5107 5364 6040 5390
rect 3340 5356 6040 5364
rect 6074 5356 6108 5390
rect 6142 5356 6176 5390
rect 6210 5356 6244 5390
rect 6278 5356 6312 5390
rect 6346 5356 6380 5390
rect 6414 5356 6448 5390
rect 6482 5356 6516 5390
rect 6550 5356 6584 5390
rect 6618 5356 6652 5390
rect 6686 5356 6720 5390
rect 6754 5375 6781 5390
rect 6754 5356 6825 5375
rect 3340 5328 5155 5356
rect 3340 5294 3373 5328
rect 3407 5294 3441 5328
rect 3475 5294 3509 5328
rect 3543 5294 3577 5328
rect 3611 5294 3645 5328
rect 3679 5294 3713 5328
rect 3747 5294 3781 5328
rect 3815 5294 3849 5328
rect 3883 5294 3917 5328
rect 3951 5294 3985 5328
rect 4019 5294 4053 5328
rect 4087 5294 4121 5328
rect 4155 5294 4189 5328
rect 4223 5294 4257 5328
rect 4291 5294 4325 5328
rect 4359 5294 4393 5328
rect 4427 5294 4461 5328
rect 4495 5294 4529 5328
rect 4563 5294 4597 5328
rect 4631 5294 4665 5328
rect 4699 5294 4733 5328
rect 4767 5294 4801 5328
rect 4835 5294 4869 5328
rect 4903 5294 4937 5328
rect 4971 5294 5005 5328
rect 5039 5294 5073 5328
rect 5107 5322 5155 5328
rect 5189 5322 5223 5356
rect 5257 5322 5291 5356
rect 5325 5322 5359 5356
rect 5393 5322 5427 5356
rect 5461 5322 5495 5356
rect 5529 5322 5563 5356
rect 5597 5322 5631 5356
rect 5665 5322 5699 5356
rect 5733 5322 5767 5356
rect 5801 5322 5835 5356
rect 5869 5322 5903 5356
rect 5937 5322 5971 5356
rect 6005 5341 6825 5356
rect 6859 5341 6893 5375
rect 6927 5341 6961 5375
rect 6995 5341 7029 5375
rect 7063 5341 7097 5375
rect 7131 5341 7165 5375
rect 7199 5341 7233 5375
rect 7267 5341 7301 5375
rect 7335 5341 7369 5375
rect 7403 5341 7437 5375
rect 7471 5341 7505 5375
rect 7539 5341 7573 5375
rect 7607 5341 7641 5375
rect 7675 5341 7709 5375
rect 7743 5341 7777 5375
rect 7811 5341 7845 5375
rect 7879 5341 7913 5375
rect 7947 5341 7981 5375
rect 8015 5341 8049 5375
rect 8083 5341 8117 5375
rect 8151 5341 8185 5375
rect 8219 5341 8253 5375
rect 8287 5341 8321 5375
rect 8355 5341 8389 5375
rect 8423 5341 8457 5375
rect 8491 5341 8525 5375
rect 8559 5341 8593 5375
rect 8627 5341 8661 5375
rect 8695 5341 8729 5375
rect 8763 5341 8797 5375
rect 8831 5341 8865 5375
rect 8899 5341 8933 5375
rect 8967 5341 9001 5375
rect 9035 5341 9069 5375
rect 9103 5341 9137 5375
rect 9171 5341 9205 5375
rect 9239 5341 9273 5375
rect 9307 5341 9341 5375
rect 9375 5341 9409 5375
rect 9443 5341 9477 5375
rect 9511 5341 9545 5375
rect 9579 5341 9613 5375
rect 9647 5341 9681 5375
rect 9715 5341 9749 5375
rect 9783 5341 9817 5375
rect 9851 5341 9886 5375
rect 9920 5341 9955 5375
rect 9989 5341 10024 5375
rect 10058 5341 10093 5375
rect 10127 5341 10162 5375
rect 10196 5341 10231 5375
rect 10265 5341 10300 5375
rect 10334 5341 10369 5375
rect 10403 5341 10438 5375
rect 10472 5341 10507 5375
rect 10541 5341 10576 5375
rect 10610 5341 10645 5375
rect 10679 5341 10714 5375
rect 10748 5341 10783 5375
rect 10817 5341 10852 5375
rect 10886 5341 10921 5375
rect 10955 5341 10990 5375
rect 11024 5341 11059 5375
rect 11093 5341 11128 5375
rect 11162 5341 11197 5375
rect 11231 5341 11266 5375
rect 11300 5341 11335 5375
rect 11369 5341 11404 5375
rect 11438 5341 11473 5375
rect 11507 5341 11542 5375
rect 11576 5341 11611 5375
rect 11645 5341 11680 5375
rect 11714 5341 11749 5375
rect 11783 5341 11818 5375
rect 11852 5341 11887 5375
rect 11921 5341 11956 5375
rect 11990 5341 12025 5375
rect 12059 5341 12094 5375
rect 12128 5341 12163 5375
rect 12197 5341 12232 5375
rect 12266 5341 12301 5375
rect 12335 5341 12370 5375
rect 12404 5341 12439 5375
rect 12473 5341 12508 5375
rect 12542 5341 12577 5375
rect 12611 5341 12646 5375
rect 12680 5341 12715 5375
rect 12749 5341 12784 5375
rect 12818 5341 12853 5375
rect 12887 5341 12922 5375
rect 12956 5341 12991 5375
rect 13025 5341 13060 5375
rect 13094 5341 13129 5375
rect 13163 5341 13197 5375
rect 6005 5322 6781 5341
rect 5107 5321 6781 5322
rect 5107 5294 6040 5321
rect 3340 5287 6040 5294
rect 6074 5287 6108 5321
rect 6142 5287 6176 5321
rect 6210 5287 6244 5321
rect 6278 5287 6312 5321
rect 6346 5287 6380 5321
rect 6414 5287 6448 5321
rect 6482 5287 6516 5321
rect 6550 5287 6584 5321
rect 6618 5287 6652 5321
rect 6686 5287 6720 5321
rect 6754 5287 6781 5321
rect 3340 5281 6781 5287
rect 3340 5257 5155 5281
rect 3340 5223 3373 5257
rect 3407 5223 3441 5257
rect 3475 5223 3509 5257
rect 3543 5223 3577 5257
rect 3611 5223 3645 5257
rect 3679 5223 3713 5257
rect 3747 5223 3781 5257
rect 3815 5223 3849 5257
rect 3883 5223 3917 5257
rect 3951 5223 3985 5257
rect 4019 5223 4053 5257
rect 4087 5223 4121 5257
rect 4155 5223 4189 5257
rect 4223 5223 4257 5257
rect 4291 5223 4325 5257
rect 4359 5223 4393 5257
rect 4427 5223 4461 5257
rect 4495 5223 4529 5257
rect 4563 5223 4597 5257
rect 4631 5223 4665 5257
rect 4699 5223 4733 5257
rect 4767 5223 4801 5257
rect 4835 5223 4869 5257
rect 4903 5223 4937 5257
rect 4971 5223 5005 5257
rect 5039 5223 5073 5257
rect 5107 5247 5155 5257
rect 5189 5247 5223 5281
rect 5257 5247 5291 5281
rect 5325 5247 5359 5281
rect 5393 5247 5427 5281
rect 5461 5247 5495 5281
rect 5529 5247 5563 5281
rect 5597 5247 5631 5281
rect 5665 5247 5699 5281
rect 5733 5247 5767 5281
rect 5801 5247 5835 5281
rect 5869 5247 5903 5281
rect 5937 5247 5971 5281
rect 6005 5251 6781 5281
rect 6005 5247 6040 5251
rect 5107 5223 6040 5247
rect 3340 5217 6040 5223
rect 6074 5217 6108 5251
rect 6142 5217 6176 5251
rect 6210 5217 6244 5251
rect 6278 5217 6312 5251
rect 6346 5217 6380 5251
rect 6414 5217 6448 5251
rect 6482 5217 6516 5251
rect 6550 5217 6584 5251
rect 6618 5217 6652 5251
rect 6686 5217 6720 5251
rect 6754 5217 6781 5251
rect 3340 5206 6781 5217
rect 3340 5186 5155 5206
rect 3340 5152 3373 5186
rect 3407 5152 3441 5186
rect 3475 5152 3509 5186
rect 3543 5152 3577 5186
rect 3611 5152 3645 5186
rect 3679 5152 3713 5186
rect 3747 5152 3781 5186
rect 3815 5152 3849 5186
rect 3883 5152 3917 5186
rect 3951 5152 3985 5186
rect 4019 5152 4053 5186
rect 4087 5152 4121 5186
rect 4155 5152 4189 5186
rect 4223 5152 4257 5186
rect 4291 5152 4325 5186
rect 4359 5152 4393 5186
rect 4427 5152 4461 5186
rect 4495 5152 4529 5186
rect 4563 5152 4597 5186
rect 4631 5152 4665 5186
rect 4699 5152 4733 5186
rect 4767 5152 4801 5186
rect 4835 5152 4869 5186
rect 4903 5152 4937 5186
rect 4971 5152 5005 5186
rect 5039 5152 5073 5186
rect 5107 5172 5155 5186
rect 5189 5172 5223 5206
rect 5257 5172 5291 5206
rect 5325 5172 5359 5206
rect 5393 5172 5427 5206
rect 5461 5172 5495 5206
rect 5529 5172 5563 5206
rect 5597 5172 5631 5206
rect 5665 5172 5699 5206
rect 5733 5172 5767 5206
rect 5801 5172 5835 5206
rect 5869 5172 5903 5206
rect 5937 5172 5971 5206
rect 6005 5181 6781 5206
rect 6005 5172 6040 5181
rect 5107 5152 6040 5172
rect 3340 5147 6040 5152
rect 6074 5147 6108 5181
rect 6142 5147 6176 5181
rect 6210 5147 6244 5181
rect 6278 5147 6312 5181
rect 6346 5147 6380 5181
rect 6414 5147 6448 5181
rect 6482 5147 6516 5181
rect 6550 5147 6584 5181
rect 6618 5147 6652 5181
rect 6686 5147 6720 5181
rect 6754 5147 6781 5181
rect 3340 5131 6781 5147
rect 3340 5115 5155 5131
rect 3340 5081 3373 5115
rect 3407 5081 3441 5115
rect 3475 5081 3509 5115
rect 3543 5081 3577 5115
rect 3611 5081 3645 5115
rect 3679 5081 3713 5115
rect 3747 5081 3781 5115
rect 3815 5081 3849 5115
rect 3883 5081 3917 5115
rect 3951 5081 3985 5115
rect 4019 5081 4053 5115
rect 4087 5081 4121 5115
rect 4155 5081 4189 5115
rect 4223 5081 4257 5115
rect 4291 5081 4325 5115
rect 4359 5081 4393 5115
rect 4427 5081 4461 5115
rect 4495 5081 4529 5115
rect 4563 5081 4597 5115
rect 4631 5081 4665 5115
rect 4699 5081 4733 5115
rect 4767 5081 4801 5115
rect 4835 5081 4869 5115
rect 4903 5081 4937 5115
rect 4971 5081 5005 5115
rect 5039 5081 5073 5115
rect 5107 5097 5155 5115
rect 5189 5097 5223 5131
rect 5257 5097 5291 5131
rect 5325 5097 5359 5131
rect 5393 5097 5427 5131
rect 5461 5097 5495 5131
rect 5529 5097 5563 5131
rect 5597 5097 5631 5131
rect 5665 5097 5699 5131
rect 5733 5097 5767 5131
rect 5801 5097 5835 5131
rect 5869 5097 5903 5131
rect 5937 5097 5971 5131
rect 6005 5111 6781 5131
rect 6852 5244 6886 5251
rect 6966 5245 7005 5279
rect 7039 5245 7078 5279
rect 7112 5245 7151 5279
rect 7185 5245 7224 5279
rect 7258 5245 7297 5279
rect 7331 5245 7370 5279
rect 7404 5245 7443 5279
rect 7477 5245 7516 5279
rect 7550 5245 7589 5279
rect 7623 5245 7662 5279
rect 7696 5245 7735 5279
rect 7769 5245 7808 5279
rect 7842 5245 7881 5279
rect 7915 5245 7954 5279
rect 7988 5245 8027 5279
rect 8061 5245 8100 5279
rect 8134 5245 8173 5279
rect 8207 5245 8246 5279
rect 8280 5245 8319 5279
rect 8353 5245 8392 5279
rect 8426 5245 8465 5279
rect 8499 5245 8538 5279
rect 8572 5245 8611 5279
rect 8645 5245 8684 5279
rect 8718 5245 8757 5279
rect 8791 5245 8830 5279
rect 8864 5245 8903 5279
rect 8937 5245 8976 5279
rect 9010 5245 9049 5279
rect 9083 5245 9122 5279
rect 9156 5245 9195 5279
rect 9229 5245 9268 5279
rect 9302 5245 9341 5279
rect 9375 5245 9414 5279
rect 9448 5245 9486 5279
rect 9520 5245 9558 5279
rect 9592 5245 9630 5279
rect 9664 5245 9702 5279
rect 9736 5245 9774 5279
rect 9808 5245 9846 5279
rect 10165 5245 10203 5279
rect 10237 5245 10275 5279
rect 10309 5245 10347 5279
rect 10381 5245 10419 5279
rect 10453 5245 10491 5279
rect 10525 5245 10563 5279
rect 10597 5245 10635 5279
rect 10669 5245 10707 5279
rect 10741 5245 10779 5279
rect 10813 5245 10852 5279
rect 10886 5245 10925 5279
rect 10959 5245 10998 5279
rect 11032 5245 11071 5279
rect 11105 5245 11144 5279
rect 11178 5245 11217 5279
rect 11251 5245 11290 5279
rect 11324 5245 11363 5279
rect 11397 5245 11436 5279
rect 11470 5245 11509 5279
rect 11543 5245 11582 5279
rect 11616 5245 11655 5279
rect 11689 5245 11728 5279
rect 11762 5245 11801 5279
rect 11835 5245 11874 5279
rect 11908 5245 11947 5279
rect 11981 5245 12020 5279
rect 12054 5245 12093 5279
rect 12127 5245 12166 5279
rect 12200 5245 12239 5279
rect 12273 5245 12312 5279
rect 12346 5245 12385 5279
rect 12419 5245 12458 5279
rect 12492 5245 12531 5279
rect 12565 5245 12604 5279
rect 12638 5245 12677 5279
rect 12711 5245 12750 5279
rect 12784 5245 12823 5279
rect 12857 5245 12896 5279
rect 12930 5245 12969 5279
rect 13003 5245 13042 5279
rect 6852 5172 6886 5201
rect 13156 5235 13159 5251
rect 13122 5201 13125 5218
rect 13122 5180 13159 5201
rect 13156 5167 13159 5180
rect 6852 5117 6886 5133
rect 6005 5097 6040 5111
rect 5107 5081 6040 5097
rect 3340 5077 6040 5081
rect 6074 5077 6108 5111
rect 6142 5077 6176 5111
rect 6210 5077 6244 5111
rect 6278 5077 6312 5111
rect 6346 5077 6380 5111
rect 6414 5077 6448 5111
rect 6482 5077 6516 5111
rect 6550 5077 6584 5111
rect 6618 5077 6652 5111
rect 6686 5077 6720 5111
rect 6754 5077 6781 5111
rect 6966 5089 7006 5123
rect 7040 5089 7080 5123
rect 7114 5089 7154 5123
rect 7188 5089 7228 5123
rect 7262 5089 7302 5123
rect 7336 5089 7376 5123
rect 7410 5089 7450 5123
rect 7484 5089 7524 5123
rect 7558 5089 7597 5123
rect 7631 5089 7670 5123
rect 7704 5089 7743 5123
rect 7777 5089 7816 5123
rect 7850 5089 7889 5123
rect 7923 5089 7962 5123
rect 7996 5089 8035 5123
rect 8069 5089 8108 5123
rect 8142 5089 8181 5123
rect 8215 5089 8254 5123
rect 8288 5089 8327 5123
rect 8361 5089 8400 5123
rect 8434 5089 8473 5123
rect 8507 5089 8546 5123
rect 8580 5089 8619 5123
rect 8653 5089 8692 5123
rect 8726 5089 8765 5123
rect 8799 5089 8838 5123
rect 8872 5089 8911 5123
rect 8945 5089 8984 5123
rect 9018 5089 9057 5123
rect 9091 5089 9130 5123
rect 9164 5089 9203 5123
rect 9237 5089 9276 5123
rect 9310 5089 9349 5123
rect 9383 5089 9422 5123
rect 9456 5089 9495 5123
rect 9529 5089 9568 5123
rect 9602 5089 9641 5123
rect 9675 5089 9714 5123
rect 9748 5089 9787 5123
rect 10230 5089 10268 5123
rect 10302 5089 10341 5123
rect 10375 5089 10414 5123
rect 10448 5089 10487 5123
rect 10521 5089 10560 5123
rect 10594 5089 10633 5123
rect 10667 5089 10706 5123
rect 10740 5089 10779 5123
rect 10813 5089 10852 5123
rect 10886 5089 10925 5123
rect 10959 5089 10998 5123
rect 11032 5089 11071 5123
rect 11105 5089 11144 5123
rect 11178 5089 11217 5123
rect 11251 5089 11290 5123
rect 11324 5089 11363 5123
rect 11397 5089 11436 5123
rect 11470 5089 11509 5123
rect 11543 5089 11582 5123
rect 11616 5089 11655 5123
rect 11689 5089 11728 5123
rect 11762 5089 11801 5123
rect 11835 5089 11874 5123
rect 11908 5089 11947 5123
rect 11981 5089 12020 5123
rect 12054 5089 12093 5123
rect 12127 5089 12166 5123
rect 12200 5089 12239 5123
rect 12273 5089 12312 5123
rect 12346 5089 12385 5123
rect 12419 5089 12458 5123
rect 12492 5089 12531 5123
rect 12565 5089 12604 5123
rect 12638 5089 12677 5123
rect 12711 5089 12750 5123
rect 12784 5089 12823 5123
rect 12857 5089 12896 5123
rect 12930 5089 12969 5123
rect 13003 5089 13042 5123
rect 13125 5117 13159 5133
rect 3340 5056 6781 5077
rect 3340 5044 5155 5056
rect 3340 5010 3373 5044
rect 3407 5010 3441 5044
rect 3475 5010 3509 5044
rect 3543 5010 3577 5044
rect 3611 5010 3645 5044
rect 3679 5010 3713 5044
rect 3747 5010 3781 5044
rect 3815 5010 3849 5044
rect 3883 5010 3917 5044
rect 3951 5010 3985 5044
rect 4019 5010 4053 5044
rect 4087 5010 4121 5044
rect 4155 5010 4189 5044
rect 4223 5010 4257 5044
rect 4291 5010 4325 5044
rect 4359 5010 4393 5044
rect 4427 5010 4461 5044
rect 4495 5010 4529 5044
rect 4563 5010 4597 5044
rect 4631 5010 4665 5044
rect 4699 5010 4733 5044
rect 4767 5010 4801 5044
rect 4835 5010 4869 5044
rect 4903 5010 4937 5044
rect 4971 5010 5005 5044
rect 5039 5010 5073 5044
rect 5107 5022 5155 5044
rect 5189 5022 5223 5056
rect 5257 5022 5291 5056
rect 5325 5022 5359 5056
rect 5393 5022 5427 5056
rect 5461 5022 5495 5056
rect 5529 5022 5563 5056
rect 5597 5022 5631 5056
rect 5665 5022 5699 5056
rect 5733 5022 5767 5056
rect 5801 5022 5835 5056
rect 5869 5022 5903 5056
rect 5937 5022 5971 5056
rect 6005 5041 6781 5056
rect 6005 5022 6040 5041
rect 5107 5010 6040 5022
rect 3340 5007 6040 5010
rect 6074 5007 6108 5041
rect 6142 5007 6176 5041
rect 6210 5007 6244 5041
rect 6278 5007 6312 5041
rect 6346 5007 6380 5041
rect 6414 5007 6448 5041
rect 6482 5007 6516 5041
rect 6550 5007 6584 5041
rect 6618 5007 6652 5041
rect 6686 5007 6720 5041
rect 6754 5007 6781 5041
rect 3340 4985 6781 5007
rect 3340 4981 6829 4985
rect 3340 4973 5155 4981
rect 3340 4939 3373 4973
rect 3407 4939 3441 4973
rect 3475 4939 3509 4973
rect 3543 4939 3577 4973
rect 3611 4939 3645 4973
rect 3679 4939 3713 4973
rect 3747 4939 3781 4973
rect 3815 4939 3849 4973
rect 3883 4939 3917 4973
rect 3951 4939 3985 4973
rect 4019 4939 4053 4973
rect 4087 4939 4121 4973
rect 4155 4939 4189 4973
rect 4223 4939 4257 4973
rect 4291 4939 4325 4973
rect 4359 4939 4393 4973
rect 4427 4939 4461 4973
rect 4495 4939 4529 4973
rect 4563 4939 4597 4973
rect 4631 4939 4665 4973
rect 4699 4939 4733 4973
rect 4767 4939 4801 4973
rect 4835 4939 4869 4973
rect 4903 4939 4937 4973
rect 4971 4939 5005 4973
rect 5039 4939 5073 4973
rect 5107 4947 5155 4973
rect 5189 4947 5223 4981
rect 5257 4947 5291 4981
rect 5325 4947 5359 4981
rect 5393 4947 5427 4981
rect 5461 4947 5495 4981
rect 5529 4947 5563 4981
rect 5597 4947 5631 4981
rect 5665 4947 5699 4981
rect 5733 4947 5767 4981
rect 5801 4947 5835 4981
rect 5869 4947 5903 4981
rect 5937 4947 5971 4981
rect 6005 4971 6829 4981
rect 6005 4947 6040 4971
rect 5107 4939 6040 4947
rect 3340 4937 6040 4939
rect 6074 4937 6108 4971
rect 6142 4937 6176 4971
rect 6210 4937 6244 4971
rect 6278 4937 6312 4971
rect 6346 4937 6380 4971
rect 6414 4937 6448 4971
rect 6482 4937 6516 4971
rect 6550 4937 6584 4971
rect 6618 4937 6652 4971
rect 6686 4937 6720 4971
rect 6754 4951 6829 4971
rect 6863 4951 6898 4985
rect 6932 4951 6967 4985
rect 7001 4951 7036 4985
rect 7070 4951 7105 4985
rect 7139 4951 7174 4985
rect 7208 4951 7243 4985
rect 7277 4951 7312 4985
rect 7346 4951 7381 4985
rect 7415 4951 7450 4985
rect 7484 4951 7519 4985
rect 7553 4951 7588 4985
rect 7622 4951 7657 4985
rect 7691 4951 7726 4985
rect 7760 4951 7795 4985
rect 7829 4951 7864 4985
rect 7898 4951 7933 4985
rect 7967 4951 8002 4985
rect 8036 4951 8071 4985
rect 8105 4951 8140 4985
rect 8174 4951 8209 4985
rect 8243 4951 8278 4985
rect 8312 4951 8347 4985
rect 8381 4951 8416 4985
rect 8450 4951 8485 4985
rect 8519 4951 8554 4985
rect 8588 4951 8623 4985
rect 6754 4937 8623 4951
rect 3340 4917 8623 4937
rect 3340 4906 6829 4917
rect 3340 4902 5155 4906
rect 3340 4868 3373 4902
rect 3407 4868 3441 4902
rect 3475 4868 3509 4902
rect 3543 4868 3577 4902
rect 3611 4868 3645 4902
rect 3679 4868 3713 4902
rect 3747 4868 3781 4902
rect 3815 4868 3849 4902
rect 3883 4868 3917 4902
rect 3951 4868 3985 4902
rect 4019 4868 4053 4902
rect 4087 4868 4121 4902
rect 4155 4868 4189 4902
rect 4223 4868 4257 4902
rect 4291 4868 4325 4902
rect 4359 4868 4393 4902
rect 4427 4868 4461 4902
rect 4495 4868 4529 4902
rect 4563 4868 4597 4902
rect 4631 4868 4665 4902
rect 4699 4868 4733 4902
rect 4767 4868 4801 4902
rect 4835 4868 4869 4902
rect 4903 4868 4937 4902
rect 4971 4868 5005 4902
rect 5039 4868 5073 4902
rect 5107 4872 5155 4902
rect 5189 4872 5223 4906
rect 5257 4872 5291 4906
rect 5325 4872 5359 4906
rect 5393 4872 5427 4906
rect 5461 4872 5495 4906
rect 5529 4872 5563 4906
rect 5597 4872 5631 4906
rect 5665 4872 5699 4906
rect 5733 4872 5767 4906
rect 5801 4872 5835 4906
rect 5869 4872 5903 4906
rect 5937 4872 5971 4906
rect 6005 4901 6829 4906
rect 6005 4872 6040 4901
rect 5107 4868 6040 4872
rect 3340 4867 6040 4868
rect 6074 4867 6108 4901
rect 6142 4867 6176 4901
rect 6210 4867 6244 4901
rect 6278 4867 6312 4901
rect 6346 4867 6380 4901
rect 6414 4867 6448 4901
rect 6482 4867 6516 4901
rect 6550 4867 6584 4901
rect 6618 4867 6652 4901
rect 6686 4867 6720 4901
rect 6754 4883 6829 4901
rect 6863 4883 6898 4917
rect 6932 4883 6967 4917
rect 7001 4883 7036 4917
rect 7070 4883 7105 4917
rect 7139 4883 7174 4917
rect 7208 4883 7243 4917
rect 7277 4883 7312 4917
rect 7346 4883 7381 4917
rect 7415 4883 7450 4917
rect 7484 4883 7519 4917
rect 7553 4883 7588 4917
rect 7622 4883 7657 4917
rect 7691 4883 7726 4917
rect 7760 4883 7795 4917
rect 7829 4883 7864 4917
rect 7898 4883 7933 4917
rect 7967 4883 8002 4917
rect 8036 4883 8071 4917
rect 8105 4883 8140 4917
rect 8174 4883 8209 4917
rect 8243 4883 8278 4917
rect 8312 4883 8347 4917
rect 8381 4883 8416 4917
rect 8450 4883 8485 4917
rect 8519 4883 8554 4917
rect 8588 4883 8623 4917
rect 6754 4867 8623 4883
rect 3340 4849 8623 4867
rect 3340 4831 6829 4849
rect 3340 4797 3373 4831
rect 3407 4797 3441 4831
rect 3475 4797 3509 4831
rect 3543 4797 3577 4831
rect 3611 4797 3645 4831
rect 3679 4797 3713 4831
rect 3747 4797 3781 4831
rect 3815 4797 3849 4831
rect 3883 4797 3917 4831
rect 3951 4797 3985 4831
rect 4019 4797 4053 4831
rect 4087 4797 4121 4831
rect 4155 4797 4189 4831
rect 4223 4797 4257 4831
rect 4291 4797 4325 4831
rect 4359 4797 4393 4831
rect 4427 4797 4461 4831
rect 4495 4797 4529 4831
rect 4563 4797 4597 4831
rect 4631 4797 4665 4831
rect 4699 4797 4733 4831
rect 4767 4797 4801 4831
rect 4835 4797 4869 4831
rect 4903 4797 4937 4831
rect 4971 4797 5005 4831
rect 5039 4797 5073 4831
rect 5107 4797 5155 4831
rect 5189 4797 5223 4831
rect 5257 4797 5291 4831
rect 5325 4797 5359 4831
rect 5393 4797 5427 4831
rect 5461 4797 5495 4831
rect 5529 4797 5563 4831
rect 5597 4797 5631 4831
rect 5665 4797 5699 4831
rect 5733 4797 5767 4831
rect 5801 4797 5835 4831
rect 5869 4797 5903 4831
rect 5937 4797 5971 4831
rect 6005 4797 6040 4831
rect 6074 4797 6108 4831
rect 6142 4797 6176 4831
rect 6210 4797 6244 4831
rect 6278 4797 6312 4831
rect 6346 4797 6380 4831
rect 6414 4797 6448 4831
rect 6482 4797 6516 4831
rect 6550 4797 6584 4831
rect 6618 4797 6652 4831
rect 6686 4797 6720 4831
rect 6754 4815 6829 4831
rect 6863 4815 6898 4849
rect 6932 4815 6967 4849
rect 7001 4815 7036 4849
rect 7070 4815 7105 4849
rect 7139 4815 7174 4849
rect 7208 4815 7243 4849
rect 7277 4815 7312 4849
rect 7346 4815 7381 4849
rect 7415 4815 7450 4849
rect 7484 4815 7519 4849
rect 7553 4815 7588 4849
rect 7622 4815 7657 4849
rect 7691 4815 7726 4849
rect 7760 4815 7795 4849
rect 7829 4815 7864 4849
rect 7898 4815 7933 4849
rect 7967 4815 8002 4849
rect 8036 4815 8071 4849
rect 8105 4815 8140 4849
rect 8174 4815 8209 4849
rect 8243 4815 8278 4849
rect 8312 4815 8347 4849
rect 8381 4815 8416 4849
rect 8450 4815 8485 4849
rect 8519 4815 8554 4849
rect 8588 4815 8623 4849
rect 13145 4815 13197 4985
rect 6754 4798 13197 4815
rect 6754 4797 13265 4798
rect 3340 4763 13265 4797
rect 3340 4729 3374 4763
rect 3408 4731 3443 4763
rect 3477 4731 3512 4763
rect 3546 4731 3581 4763
rect 3615 4731 3650 4763
rect 3684 4731 3719 4763
rect 3753 4731 3788 4763
rect 3822 4731 3857 4763
rect 3891 4731 3926 4763
rect 3960 4731 3995 4763
rect 3408 4729 3410 4731
rect 3477 4729 3483 4731
rect 3546 4729 3556 4731
rect 3615 4729 3629 4731
rect 3684 4729 3702 4731
rect 3753 4729 3775 4731
rect 3822 4729 3848 4731
rect 3891 4729 3921 4731
rect 3960 4729 3994 4731
rect 4029 4729 4064 4763
rect 4098 4731 4133 4763
rect 4167 4731 4202 4763
rect 4236 4731 4271 4763
rect 4305 4731 4340 4763
rect 4374 4731 4409 4763
rect 4443 4731 4478 4763
rect 4512 4731 4547 4763
rect 4581 4731 4616 4763
rect 4101 4729 4133 4731
rect 4174 4729 4202 4731
rect 4247 4729 4271 4731
rect 4320 4729 4340 4731
rect 4393 4729 4409 4731
rect 4466 4729 4478 4731
rect 4539 4729 4547 4731
rect 4612 4729 4616 4731
rect 4650 4731 4685 4763
rect 4650 4729 4651 4731
rect 3340 4697 3410 4729
rect 3444 4697 3483 4729
rect 3517 4697 3556 4729
rect 3590 4697 3629 4729
rect 3663 4697 3702 4729
rect 3736 4697 3775 4729
rect 3809 4697 3848 4729
rect 3882 4697 3921 4729
rect 3955 4697 3994 4729
rect 4028 4697 4067 4729
rect 4101 4697 4140 4729
rect 4174 4697 4213 4729
rect 4247 4697 4286 4729
rect 4320 4697 4359 4729
rect 4393 4697 4432 4729
rect 4466 4697 4505 4729
rect 4539 4697 4578 4729
rect 4612 4697 4651 4729
rect 4719 4731 4754 4763
rect 4788 4731 4823 4763
rect 4857 4731 4892 4763
rect 4926 4731 4961 4763
rect 4995 4731 5030 4763
rect 5064 4731 5099 4763
rect 5133 4731 5168 4763
rect 5202 4731 5237 4763
rect 4719 4729 4724 4731
rect 4788 4729 4797 4731
rect 4857 4729 4870 4731
rect 4926 4729 4943 4731
rect 4995 4729 5016 4731
rect 5064 4729 5089 4731
rect 5133 4729 5162 4731
rect 5202 4729 5235 4731
rect 5271 4729 5306 4763
rect 5340 4731 5375 4763
rect 5409 4731 5444 4763
rect 5478 4731 5513 4763
rect 5547 4731 5582 4763
rect 5616 4731 5651 4763
rect 5685 4731 5720 4763
rect 5754 4731 5789 4763
rect 5823 4731 5858 4763
rect 5892 4731 5927 4763
rect 5961 4731 5996 4763
rect 6030 4731 6065 4763
rect 5341 4729 5375 4731
rect 5413 4729 5444 4731
rect 5485 4729 5513 4731
rect 5557 4729 5582 4731
rect 5629 4729 5651 4731
rect 5701 4729 5720 4731
rect 5773 4729 5789 4731
rect 5845 4729 5858 4731
rect 5917 4729 5927 4731
rect 5989 4729 5996 4731
rect 6061 4729 6065 4731
rect 6099 4731 6134 4763
rect 4685 4697 4724 4729
rect 4758 4697 4797 4729
rect 4831 4697 4870 4729
rect 4904 4697 4943 4729
rect 4977 4697 5016 4729
rect 5050 4697 5089 4729
rect 5123 4697 5162 4729
rect 5196 4697 5235 4729
rect 5269 4697 5307 4729
rect 5341 4697 5379 4729
rect 5413 4697 5451 4729
rect 5485 4697 5523 4729
rect 5557 4697 5595 4729
rect 5629 4697 5667 4729
rect 5701 4697 5739 4729
rect 5773 4697 5811 4729
rect 5845 4697 5883 4729
rect 5917 4697 5955 4729
rect 5989 4697 6027 4729
rect 6061 4697 6099 4729
rect 6133 4729 6134 4731
rect 6168 4731 6203 4763
rect 6237 4731 6272 4763
rect 6306 4731 6341 4763
rect 6375 4731 6410 4763
rect 6444 4731 6479 4763
rect 6513 4731 6548 4763
rect 6582 4731 6617 4763
rect 6651 4731 6686 4763
rect 6720 4731 6755 4763
rect 6789 4731 6824 4763
rect 6858 4731 6893 4763
rect 6168 4729 6171 4731
rect 6237 4729 6243 4731
rect 6306 4729 6315 4731
rect 6375 4729 6387 4731
rect 6444 4729 6459 4731
rect 6513 4729 6531 4731
rect 6582 4729 6603 4731
rect 6651 4729 6675 4731
rect 6720 4729 6747 4731
rect 6789 4729 6819 4731
rect 6858 4729 6891 4731
rect 6927 4729 6962 4763
rect 10056 4731 10092 4763
rect 10126 4731 10161 4763
rect 10195 4731 10230 4763
rect 10264 4731 10299 4763
rect 10333 4731 10368 4763
rect 10402 4731 10437 4763
rect 10471 4731 10506 4763
rect 10540 4731 10575 4763
rect 10609 4731 10644 4763
rect 10678 4731 10713 4763
rect 10747 4731 10782 4763
rect 10816 4731 10851 4763
rect 10885 4731 10920 4763
rect 10954 4731 10989 4763
rect 11023 4731 11058 4763
rect 11092 4731 11127 4763
rect 11161 4731 11196 4763
rect 11230 4731 11265 4763
rect 11299 4731 11334 4763
rect 11368 4731 11403 4763
rect 11437 4731 11472 4763
rect 11506 4731 11541 4763
rect 11575 4731 11610 4763
rect 11644 4731 11679 4763
rect 11713 4731 11748 4763
rect 11782 4731 11817 4763
rect 11851 4731 11886 4763
rect 11920 4731 11955 4763
rect 11989 4731 12024 4763
rect 12058 4731 12093 4763
rect 12127 4731 12162 4763
rect 12196 4731 12231 4763
rect 12265 4731 12300 4763
rect 12334 4731 12369 4763
rect 12403 4731 12438 4763
rect 12472 4731 12507 4763
rect 12541 4731 12576 4763
rect 12610 4731 12645 4763
rect 12679 4731 12714 4763
rect 12748 4731 12783 4763
rect 12817 4731 12852 4763
rect 12886 4731 12921 4763
rect 12955 4731 12990 4763
rect 13024 4731 13059 4763
rect 13093 4731 13128 4763
rect 13162 4731 13197 4763
rect 13231 4731 13265 4763
rect 6133 4697 6171 4729
rect 6205 4697 6243 4729
rect 6277 4697 6315 4729
rect 6349 4697 6387 4729
rect 6421 4697 6459 4729
rect 6493 4697 6531 4729
rect 6565 4697 6603 4729
rect 6637 4697 6675 4729
rect 6709 4697 6747 4729
rect 6781 4697 6819 4729
rect 6853 4697 6891 4729
rect 6925 4697 6962 4729
rect 3340 4695 6962 4697
rect 3340 4661 3408 4695
rect 3442 4661 3477 4695
rect 3511 4661 3546 4695
rect 3580 4661 3615 4695
rect 3649 4661 3684 4695
rect 3718 4661 3753 4695
rect 3787 4661 3822 4695
rect 3856 4661 3891 4695
rect 3925 4661 3960 4695
rect 3994 4661 4029 4695
rect 4063 4661 4098 4695
rect 4132 4661 4167 4695
rect 4201 4661 4236 4695
rect 4270 4661 4305 4695
rect 4339 4661 4374 4695
rect 4408 4661 4443 4695
rect 4477 4661 4512 4695
rect 4546 4661 4581 4695
rect 4615 4661 4650 4695
rect 4684 4661 4718 4695
rect 3340 4659 4718 4661
rect 3340 4657 3444 4659
rect 3374 4625 3444 4657
rect 3478 4627 3517 4659
rect 3551 4627 3590 4659
rect 3624 4627 3663 4659
rect 3697 4627 3736 4659
rect 3770 4627 3809 4659
rect 3843 4627 3882 4659
rect 3916 4627 3955 4659
rect 3989 4627 4028 4659
rect 4062 4627 4101 4659
rect 4135 4627 4174 4659
rect 4208 4627 4247 4659
rect 4281 4627 4320 4659
rect 4354 4627 4393 4659
rect 4427 4627 4466 4659
rect 4500 4627 4539 4659
rect 4573 4627 4612 4659
rect 4646 4627 4685 4659
rect 3510 4625 3517 4627
rect 3579 4625 3590 4627
rect 3648 4625 3663 4627
rect 3717 4625 3736 4627
rect 3786 4625 3809 4627
rect 3855 4625 3882 4627
rect 3924 4625 3955 4627
rect 3374 4623 3476 4625
rect 3340 4622 3476 4623
rect 3340 4613 3408 4622
rect 3340 4587 3372 4613
rect 3406 4588 3408 4613
rect 3442 4593 3476 4622
rect 3510 4593 3545 4625
rect 3579 4593 3614 4625
rect 3648 4593 3683 4625
rect 3717 4593 3752 4625
rect 3786 4593 3821 4625
rect 3855 4593 3890 4625
rect 3924 4593 3959 4625
rect 3993 4593 4028 4627
rect 4062 4593 4097 4627
rect 4135 4625 4166 4627
rect 4208 4625 4235 4627
rect 4281 4625 4304 4627
rect 4354 4625 4373 4627
rect 4427 4625 4442 4627
rect 4500 4625 4511 4627
rect 4573 4625 4580 4627
rect 4646 4625 4649 4627
rect 4131 4593 4166 4625
rect 4200 4593 4235 4625
rect 4269 4593 4304 4625
rect 4338 4593 4373 4625
rect 4407 4593 4442 4625
rect 4476 4593 4511 4625
rect 4545 4593 4580 4625
rect 4614 4593 4649 4625
rect 4683 4625 4685 4627
rect 13333 4661 13367 4696
rect 13333 4625 13367 4627
rect 4683 4593 4718 4625
rect 10056 4593 10091 4625
rect 10125 4593 10160 4625
rect 10194 4593 10229 4625
rect 10263 4593 10298 4625
rect 10332 4593 10367 4625
rect 10401 4593 10436 4625
rect 10470 4593 10505 4625
rect 10539 4593 10574 4625
rect 10608 4593 10643 4625
rect 10677 4593 10712 4625
rect 10746 4593 10781 4625
rect 10815 4593 10850 4625
rect 10884 4593 10919 4625
rect 10953 4593 10987 4625
rect 11021 4593 11055 4625
rect 11089 4593 11123 4625
rect 11157 4593 11191 4625
rect 11225 4593 11259 4625
rect 11293 4593 11327 4625
rect 11361 4593 11395 4625
rect 11429 4593 11463 4625
rect 11497 4593 11531 4625
rect 11565 4593 11599 4625
rect 11633 4593 11667 4625
rect 11701 4593 11735 4625
rect 11769 4593 11803 4625
rect 11837 4593 11871 4625
rect 11905 4593 11939 4625
rect 11973 4593 12007 4625
rect 12041 4593 12075 4625
rect 12109 4593 12143 4625
rect 12177 4593 12211 4625
rect 12245 4593 12279 4625
rect 12313 4593 12347 4625
rect 12381 4593 12415 4625
rect 12449 4593 12483 4625
rect 12517 4593 12551 4625
rect 12585 4593 12619 4625
rect 12653 4593 12687 4625
rect 12721 4593 12755 4625
rect 12789 4593 12823 4625
rect 12857 4593 12891 4625
rect 12925 4593 12959 4625
rect 12993 4593 13027 4625
rect 13061 4593 13095 4625
rect 13129 4593 13163 4625
rect 13197 4593 13231 4625
rect 13265 4593 13367 4625
rect 3442 4588 3510 4593
rect 3406 4582 3510 4588
rect 3406 4579 3444 4582
rect 3374 4553 3444 4579
rect 3478 4557 3510 4582
rect 3340 4549 3444 4553
rect 3340 4537 3408 4549
rect 3340 4517 3372 4537
rect 3406 4515 3408 4537
rect 3442 4548 3444 4549
rect 3442 4523 3476 4548
rect 3442 4515 3510 4523
rect 3406 4505 3510 4515
rect 3406 4503 3444 4505
rect 3374 4483 3444 4503
rect 3478 4487 3510 4505
rect 3340 4476 3444 4483
rect 3340 4461 3408 4476
rect 3340 4447 3372 4461
rect 3406 4442 3408 4461
rect 3442 4471 3444 4476
rect 3442 4453 3476 4471
rect 3442 4442 3510 4453
rect 3406 4428 3510 4442
rect 3406 4427 3444 4428
rect 3374 4413 3444 4427
rect 3478 4417 3510 4428
rect 3340 4403 3444 4413
rect 3340 4384 3408 4403
rect 3340 4377 3372 4384
rect 3406 4369 3408 4384
rect 3442 4394 3444 4403
rect 3442 4383 3476 4394
rect 3442 4369 3510 4383
rect 3406 4351 3510 4369
rect 3406 4350 3444 4351
rect 3374 4343 3444 4350
rect 3478 4347 3510 4351
rect 3340 4330 3444 4343
rect 3340 4307 3408 4330
rect 3406 4296 3408 4307
rect 3442 4317 3444 4330
rect 3442 4313 3476 4317
rect 3442 4296 3510 4313
rect 3406 4277 3510 4296
rect 3406 4274 3476 4277
rect 3406 4273 3444 4274
rect 3340 4256 3444 4273
rect 3340 4237 3408 4256
rect 3374 4230 3408 4237
rect 3406 4222 3408 4230
rect 3442 4240 3444 4256
rect 3478 4240 3510 4243
rect 3442 4222 3510 4240
rect 3406 4207 3510 4222
rect 3340 4196 3372 4203
rect 3406 4197 3476 4207
rect 3406 4196 3444 4197
rect 3340 4182 3444 4196
rect 3340 4167 3408 4182
rect 3374 4153 3408 4167
rect 3406 4148 3408 4153
rect 3442 4163 3444 4182
rect 18309 4185 18366 4602
rect 3478 4163 3510 4173
rect 3442 4148 3510 4163
rect 3406 4136 3510 4148
rect 3340 4119 3372 4133
rect 3406 4120 3476 4136
rect 3406 4119 3444 4120
rect 3340 4108 3444 4119
rect 3340 4096 3408 4108
rect 3374 4076 3408 4096
rect 3406 4074 3408 4076
rect 3442 4086 3444 4108
rect 3478 4086 3510 4102
rect 3442 4074 3510 4086
rect 3406 4065 3510 4074
rect 16111 4104 16145 4142
rect 16287 4104 16321 4142
rect 16463 4104 16497 4142
rect 16639 4104 16673 4142
rect 16837 4104 16871 4142
rect 18309 4124 18516 4185
rect 3340 4042 3372 4062
rect 3406 4043 3476 4065
rect 3406 4042 3444 4043
rect 3340 4034 3444 4042
rect 3340 4025 3408 4034
rect 3374 4000 3408 4025
rect 3442 4009 3444 4034
rect 3478 4009 3510 4031
rect 3442 4000 3510 4009
rect 3374 3999 3510 4000
rect 3406 3994 3510 3999
rect 3340 3965 3372 3991
rect 3406 3966 3476 3994
rect 3406 3965 3444 3966
rect 3340 3960 3444 3965
rect 3340 3954 3408 3960
rect -25 3920 -1 3954
rect 33 3922 68 3954
rect 102 3922 137 3954
rect 171 3922 206 3954
rect 240 3922 275 3954
rect 309 3922 344 3954
rect 378 3922 413 3954
rect 447 3922 482 3954
rect 516 3922 551 3954
rect 585 3922 620 3954
rect 3374 3926 3408 3954
rect 3442 3932 3444 3960
rect 3478 3932 3510 3960
rect 3442 3926 3510 3932
rect 3374 3923 3510 3926
rect 3374 3922 3476 3923
rect 33 3920 35 3922
rect 102 3920 108 3922
rect 171 3920 181 3922
rect 240 3920 254 3922
rect 309 3920 327 3922
rect 378 3920 400 3922
rect 447 3920 473 3922
rect 516 3920 546 3922
rect 585 3920 619 3922
rect -25 3888 35 3920
rect 69 3888 108 3920
rect 142 3888 181 3920
rect 215 3888 254 3920
rect 288 3888 327 3920
rect 361 3888 400 3920
rect 434 3888 473 3920
rect 507 3888 546 3920
rect 580 3888 619 3920
rect 3406 3889 3476 3922
rect 3406 3888 3510 3889
rect -25 3886 620 3888
rect 3374 3886 3444 3888
rect -25 3852 -1 3886
rect 33 3852 68 3886
rect 102 3852 137 3886
rect 171 3852 206 3886
rect 240 3852 275 3886
rect 309 3852 344 3886
rect 378 3852 413 3886
rect 447 3852 482 3886
rect 516 3852 551 3886
rect 585 3852 620 3886
rect 3442 3854 3444 3886
rect 3478 3854 3510 3888
rect 3442 3852 3510 3854
rect -25 3850 2966 3852
rect -25 3818 35 3850
rect 69 3818 109 3850
rect 143 3818 183 3850
rect 217 3818 257 3850
rect 291 3818 331 3850
rect 365 3818 405 3850
rect 439 3818 479 3850
rect 513 3818 553 3850
rect 587 3818 627 3850
rect 661 3818 701 3850
rect 735 3818 775 3850
rect 809 3818 849 3850
rect 883 3818 923 3850
rect 957 3818 996 3850
rect 1030 3818 1069 3850
rect -25 3784 -1 3818
rect 33 3816 35 3818
rect 102 3816 109 3818
rect 171 3816 183 3818
rect 240 3816 257 3818
rect 309 3816 331 3818
rect 378 3816 405 3818
rect 447 3816 479 3818
rect 33 3784 68 3816
rect 102 3784 137 3816
rect 171 3784 206 3816
rect 240 3784 275 3816
rect 309 3784 344 3816
rect 378 3784 413 3816
rect 447 3784 482 3816
rect 516 3784 551 3818
rect 587 3816 620 3818
rect 661 3816 689 3818
rect 735 3816 758 3818
rect 809 3816 827 3818
rect 883 3816 896 3818
rect 957 3816 965 3818
rect 1030 3816 1034 3818
rect 585 3784 620 3816
rect 654 3784 689 3816
rect 723 3784 758 3816
rect 792 3784 827 3816
rect 861 3784 896 3816
rect 930 3784 965 3816
rect 999 3784 1034 3816
rect 1068 3816 1069 3818
rect 1103 3818 1142 3850
rect 1176 3818 1215 3850
rect 1249 3818 1288 3850
rect 1322 3818 1361 3850
rect 1395 3818 1434 3850
rect 1468 3818 1507 3850
rect 1541 3818 1580 3850
rect 1614 3818 1653 3850
rect 1687 3818 1726 3850
rect 1760 3818 1799 3850
rect 1833 3818 1872 3850
rect 1906 3818 1945 3850
rect 1979 3818 2018 3850
rect 2052 3818 2091 3850
rect 2125 3818 2164 3850
rect 2198 3818 2237 3850
rect 2271 3818 2310 3850
rect 1068 3784 1103 3816
rect 1137 3816 1142 3818
rect 1206 3816 1215 3818
rect 1275 3816 1288 3818
rect 1344 3816 1361 3818
rect 1413 3816 1434 3818
rect 1482 3816 1507 3818
rect 1551 3816 1580 3818
rect 1620 3816 1653 3818
rect 1137 3784 1172 3816
rect 1206 3784 1241 3816
rect 1275 3784 1310 3816
rect 1344 3784 1379 3816
rect 1413 3784 1448 3816
rect 1482 3784 1517 3816
rect 1551 3784 1586 3816
rect 1620 3784 1655 3816
rect 1689 3784 1724 3818
rect 1760 3816 1793 3818
rect 1833 3816 1862 3818
rect 1906 3816 1931 3818
rect 1979 3816 2000 3818
rect 2052 3816 2069 3818
rect 2125 3816 2138 3818
rect 2198 3816 2207 3818
rect 2271 3816 2276 3818
rect 1758 3784 1793 3816
rect 1827 3784 1862 3816
rect 1896 3784 1931 3816
rect 1965 3784 2000 3816
rect 2034 3784 2069 3816
rect 2103 3784 2138 3816
rect 2172 3784 2207 3816
rect 2241 3784 2276 3816
rect 2344 3818 2383 3850
rect 2417 3818 2456 3850
rect 2490 3818 2529 3850
rect 2563 3818 2602 3850
rect 2636 3818 2675 3850
rect 2709 3818 2748 3850
rect 2782 3818 2821 3850
rect 2855 3818 2894 3850
rect 2928 3818 2966 3850
rect 2344 3816 2345 3818
rect 2310 3784 2345 3816
rect 2379 3816 2383 3818
rect 2448 3816 2456 3818
rect 2517 3816 2529 3818
rect 2586 3816 2602 3818
rect 2655 3816 2675 3818
rect 2724 3816 2748 3818
rect 2793 3816 2821 3818
rect 2862 3816 2894 3818
rect 2379 3784 2414 3816
rect 2448 3784 2483 3816
rect 2517 3784 2552 3816
rect 2586 3784 2621 3816
rect 2655 3784 2690 3816
rect 2724 3784 2759 3816
rect 2793 3784 2828 3816
rect 2862 3784 2897 3816
rect 2931 3784 2966 3818
rect 3408 3818 3476 3852
rect 3408 3784 3510 3818
rect 16924 3646 16958 3684
rect 18451 3590 18516 4124
rect 18367 3390 18516 3590
rect 18451 3137 18516 3390
rect 13034 3103 13425 3137
rect 13459 3103 13498 3137
rect 13532 3103 13571 3137
rect 13605 3103 13644 3137
rect 13678 3103 13717 3137
rect 13751 3103 13790 3137
rect 13824 3103 13863 3137
rect 13897 3103 13936 3137
rect 13970 3103 14009 3137
rect 14043 3103 14082 3137
rect 14116 3103 14155 3137
rect 14189 3103 14228 3137
rect 14262 3103 14301 3137
rect 14335 3103 14374 3137
rect 14408 3103 14447 3137
rect 14481 3103 14519 3137
rect 14553 3103 14591 3137
rect 14625 3103 14663 3137
rect 14697 3103 14735 3137
rect 14769 3103 14807 3137
rect 14841 3103 14879 3137
rect 14913 3103 14951 3137
rect 14985 3103 15023 3137
rect 15057 3103 15095 3137
rect 15129 3103 15167 3137
rect 15201 3103 15239 3137
rect 15273 3103 15311 3137
rect 15345 3103 15383 3137
rect 15417 3103 15455 3137
rect 15489 3103 15527 3137
rect 15561 3103 15599 3137
rect 15633 3103 15671 3137
rect 15705 3103 15743 3137
rect 15777 3103 15815 3137
rect 15849 3103 15887 3137
rect 15921 3103 15959 3137
rect 15993 3103 16031 3137
rect 16065 3103 16103 3137
rect 16137 3103 16175 3137
rect 16209 3103 16247 3137
rect 16281 3103 16319 3137
rect 16353 3103 16391 3137
rect 16425 3103 16463 3137
rect 16497 3103 16535 3137
rect 16569 3103 16607 3137
rect 16641 3103 16679 3137
rect 16713 3103 16751 3137
rect 16785 3103 16823 3137
rect 16857 3103 16895 3137
rect 16929 3103 16967 3137
rect 17001 3103 17039 3137
rect 17073 3103 17111 3137
rect 17145 3103 17183 3137
rect 17217 3103 17255 3137
rect 17289 3103 17327 3137
rect 17361 3103 17399 3137
rect 17433 3103 17471 3137
rect 17505 3103 17543 3137
rect 17577 3103 17615 3137
rect 17649 3103 17687 3137
rect 17721 3103 17759 3137
rect 17793 3103 17831 3137
rect 17865 3103 17903 3137
rect 17937 3103 17975 3137
rect 18009 3103 18047 3137
rect 18081 3103 18119 3137
rect 18153 3103 18191 3137
rect 18225 3103 18263 3137
rect 18297 3103 18335 3137
rect 18369 3103 18407 3137
rect 18441 3103 18479 3137
rect 18513 3103 18551 3137
rect 18585 3103 18623 3137
rect 18657 3103 18695 3137
rect 18729 3103 18767 3137
rect 18801 3103 18839 3137
rect 18873 3103 18911 3137
rect 18945 3103 18983 3137
rect 19017 3103 19127 3137
rect 13034 3099 19127 3103
rect 13034 3065 19093 3099
rect 13034 3023 19127 3065
rect 13034 3013 19093 3023
rect 13034 2979 13058 3013
rect 13092 2979 13127 3013
rect 13161 2979 13196 3013
rect 13230 2979 13265 3013
rect 13299 2979 13334 3013
rect 13368 2979 13403 3013
rect 13437 2979 13472 3013
rect 13506 2979 13541 3013
rect 13575 2979 13610 3013
rect 13644 2979 13679 3013
rect 13713 2979 13748 3013
rect 13782 2979 13817 3013
rect 13851 2979 13886 3013
rect 13920 2979 13955 3013
rect 13989 2979 14024 3013
rect 14058 2979 14093 3013
rect 14127 2979 14162 3013
rect 14196 2979 14231 3013
rect 14265 2979 14299 3013
rect 14333 2979 14367 3013
rect 14401 2979 14435 3013
rect 14469 2979 14503 3013
rect 14537 2979 14571 3013
rect 14605 2979 14639 3013
rect 14673 2979 14707 3013
rect 14741 2979 14775 3013
rect 14809 2979 14843 3013
rect 14877 2979 14911 3013
rect 14945 2979 14979 3013
rect 15013 2979 15047 3013
rect 15081 2979 15115 3013
rect 15149 2979 15183 3013
rect 15217 2979 15251 3013
rect 15285 2979 15319 3013
rect 15353 2979 15387 3013
rect 15421 2979 15455 3013
rect 15489 2979 15523 3013
rect 15557 2979 15591 3013
rect 15625 2979 15659 3013
rect 15693 2979 15727 3013
rect 15761 2979 15795 3013
rect 15829 2979 15863 3013
rect 15897 2979 15931 3013
rect 15965 2979 15999 3013
rect 16033 2979 16067 3013
rect 16101 2979 16135 3013
rect 16169 2979 16203 3013
rect 16237 2979 16271 3013
rect 16305 2979 16339 3013
rect 16373 2979 16407 3013
rect 16441 2979 16475 3013
rect 16509 2979 16543 3013
rect 16577 2979 16611 3013
rect 16645 2979 16679 3013
rect 16713 2979 16747 3013
rect 16781 2979 16815 3013
rect 16849 2979 16883 3013
rect 16917 2979 16951 3013
rect 16985 2979 17019 3013
rect 17053 2979 17087 3013
rect 17121 2979 17155 3013
rect 17189 2979 17223 3013
rect 17257 2979 17291 3013
rect 17325 2979 17359 3013
rect 17393 2979 17427 3013
rect 17461 2979 17495 3013
rect 17529 2979 17563 3013
rect 17597 2979 17631 3013
rect 17665 2979 17699 3013
rect 17733 2979 17767 3013
rect 17801 2979 17835 3013
rect 17869 2979 17903 3013
rect 17937 2979 17971 3013
rect 18005 2979 18039 3013
rect 19025 2989 19093 3013
rect 19127 2989 19195 3019
rect 19025 2979 19195 2989
rect 13034 2945 18067 2979
rect 19025 2945 19093 2979
rect 13034 2911 15169 2945
rect 15203 2911 15238 2945
rect 15272 2911 15307 2945
rect 15341 2911 15376 2945
rect 15410 2911 15445 2945
rect 15479 2911 15514 2945
rect 15548 2911 15583 2945
rect 15617 2911 15652 2945
rect 15686 2911 15721 2945
rect 15755 2911 15790 2945
rect 15824 2911 15859 2945
rect 15893 2911 15928 2945
rect 15962 2911 15997 2945
rect 16031 2911 16066 2945
rect 16100 2911 16135 2945
rect 16169 2911 16204 2945
rect 16238 2911 16273 2945
rect 16307 2911 16342 2945
rect 16376 2911 16411 2945
rect 16445 2911 16480 2945
rect 16514 2911 16549 2945
rect 16583 2911 16618 2945
rect 16652 2911 16687 2945
rect 16721 2911 16756 2945
rect 16790 2911 16825 2945
rect 16859 2911 16894 2945
rect 16928 2911 16963 2945
rect 16997 2911 17032 2945
rect 17066 2911 17101 2945
rect 17135 2911 17170 2945
rect 17204 2911 17239 2945
rect 17273 2911 17308 2945
rect 17342 2911 17377 2945
rect 17411 2911 17446 2945
rect 17480 2911 17515 2945
rect 17549 2911 17584 2945
rect 17618 2911 17653 2945
rect 17687 2911 17722 2945
rect 17756 2911 17791 2945
rect 17825 2911 17860 2945
rect 17894 2911 17929 2945
rect 17963 2911 17998 2945
rect 18032 2911 18067 2945
rect 13034 2877 13058 2911
rect 13092 2877 13127 2911
rect 13161 2877 13196 2911
rect 13230 2877 13265 2911
rect 13299 2877 13334 2911
rect 13368 2877 13403 2911
rect 13437 2877 13472 2911
rect 13506 2877 13541 2911
rect 13575 2877 13610 2911
rect 13644 2877 13679 2911
rect 13713 2877 13748 2911
rect 13782 2877 13817 2911
rect 13851 2877 13886 2911
rect 13920 2877 13954 2911
rect 13988 2877 14022 2911
rect 14056 2877 14090 2911
rect 14124 2877 14158 2911
rect 14192 2877 14226 2911
rect 14260 2877 14294 2911
rect 14328 2877 14362 2911
rect 14396 2877 14430 2911
rect 14464 2877 14498 2911
rect 14532 2877 14566 2911
rect 14600 2877 14634 2911
rect 14668 2877 14702 2911
rect 14736 2877 14770 2911
rect 14804 2877 14838 2911
rect 14872 2877 14906 2911
rect 14940 2877 14974 2911
rect 15008 2877 15042 2911
rect 15076 2877 18067 2911
rect 13034 2843 15169 2877
rect 15203 2843 15238 2877
rect 15272 2843 15307 2877
rect 15341 2843 15376 2877
rect 15410 2843 15445 2877
rect 15479 2843 15514 2877
rect 15548 2843 15583 2877
rect 15617 2843 15652 2877
rect 15686 2843 15721 2877
rect 15755 2843 15790 2877
rect 15824 2843 15859 2877
rect 15893 2843 15928 2877
rect 15962 2843 15997 2877
rect 16031 2843 16066 2877
rect 16100 2843 16135 2877
rect 16169 2843 16204 2877
rect 16238 2843 16273 2877
rect 16307 2843 16342 2877
rect 16376 2843 16411 2877
rect 16445 2843 16480 2877
rect 16514 2843 16549 2877
rect 16583 2843 16618 2877
rect 16652 2843 16687 2877
rect 16721 2843 16756 2877
rect 16790 2843 16825 2877
rect 16859 2843 16894 2877
rect 16928 2843 16963 2877
rect 16997 2843 17032 2877
rect 17066 2843 17101 2877
rect 17135 2843 17170 2877
rect 17204 2843 17239 2877
rect 17273 2843 17308 2877
rect 17342 2843 17377 2877
rect 17411 2843 17446 2877
rect 17480 2843 17515 2877
rect 17549 2843 17584 2877
rect 17618 2843 17653 2877
rect 17687 2843 17722 2877
rect 17756 2843 17791 2877
rect 17825 2843 17860 2877
rect 17894 2843 17929 2877
rect 17963 2843 17998 2877
rect 18032 2843 18067 2877
rect 19053 2913 19093 2945
rect 19127 2913 19195 2979
rect 19053 2910 19195 2913
rect 19053 2876 19093 2910
rect 19127 2876 19195 2910
rect 19053 2872 19195 2876
rect 19053 2843 19093 2872
rect 13034 2818 19093 2843
rect 13034 2809 13500 2818
rect 13034 2775 13058 2809
rect 13092 2775 13126 2809
rect 13160 2775 13194 2809
rect 13228 2775 13262 2809
rect 13296 2775 13330 2809
rect 13364 2775 13398 2809
rect 13432 2775 13466 2809
rect 13034 2739 13500 2775
rect 13034 2705 13058 2739
rect 13092 2705 13126 2739
rect 13160 2705 13194 2739
rect 13228 2705 13262 2739
rect 13296 2705 13330 2739
rect 13364 2705 13398 2739
rect 13432 2705 13466 2739
rect 13034 2669 13500 2705
rect 13034 2635 13058 2669
rect 13092 2635 13126 2669
rect 13160 2635 13194 2669
rect 13228 2635 13262 2669
rect 13296 2635 13330 2669
rect 13364 2635 13398 2669
rect 13432 2635 13466 2669
rect 13034 2599 13500 2635
rect 19014 2807 19093 2818
rect 19127 2807 19195 2872
rect 19014 2797 19195 2807
rect 19014 2738 19093 2797
rect 19127 2738 19195 2797
rect 19014 2722 19195 2738
rect 19014 2669 19093 2722
rect 19127 2669 19195 2722
rect 19014 2647 19195 2669
rect 19014 2601 19093 2647
rect 13034 2565 13058 2599
rect 13092 2565 13126 2599
rect 13160 2565 13194 2599
rect 13228 2565 13262 2599
rect 13296 2565 13330 2599
rect 13364 2565 13398 2599
rect 13432 2565 13466 2599
rect 13034 2529 13500 2565
rect 13034 2495 13058 2529
rect 13092 2495 13126 2529
rect 13160 2495 13194 2529
rect 13228 2495 13262 2529
rect 13296 2495 13330 2529
rect 13364 2495 13398 2529
rect 13432 2495 13466 2529
rect 13034 2460 13500 2495
rect 13034 2426 13058 2460
rect 13092 2426 13126 2460
rect 13160 2426 13194 2460
rect 13228 2426 13262 2460
rect 13296 2426 13330 2460
rect 13364 2426 13398 2460
rect 13432 2426 13466 2460
rect 19071 2600 19093 2601
rect 19127 2600 19195 2647
rect 19071 2572 19195 2600
rect 19071 2531 19093 2572
rect 19127 2531 19195 2572
rect 19071 2497 19195 2531
rect 19071 2462 19093 2497
rect 19127 2462 19195 2497
rect 19071 2438 19195 2462
rect 13034 2391 13500 2426
rect 13034 2357 13058 2391
rect 13092 2357 13126 2391
rect 13160 2357 13194 2391
rect 13228 2357 13262 2391
rect 13296 2357 13330 2391
rect 13364 2357 13398 2391
rect 13432 2357 13466 2391
rect 13034 2322 13500 2357
rect 13034 2288 13058 2322
rect 13092 2288 13126 2322
rect 13160 2288 13194 2322
rect 13228 2288 13262 2322
rect 13296 2288 13330 2322
rect 13364 2288 13398 2322
rect 13432 2288 13466 2322
rect 13034 2253 13500 2288
rect 13034 2219 13058 2253
rect 13092 2219 13126 2253
rect 13160 2219 13194 2253
rect 13228 2219 13262 2253
rect 13296 2219 13330 2253
rect 13364 2219 13398 2253
rect 13432 2219 13466 2253
rect 13034 2184 13500 2219
rect 13034 2150 13058 2184
rect 13092 2150 13126 2184
rect 13160 2150 13194 2184
rect 13228 2150 13262 2184
rect 13296 2150 13330 2184
rect 13364 2150 13398 2184
rect 13432 2150 13466 2184
rect 13034 2115 13500 2150
rect 18258 2137 18994 2249
rect 19100 2247 19193 2271
rect 19125 2213 19159 2247
rect 19100 2176 19193 2213
rect 19125 2142 19159 2176
rect 13034 2081 13058 2115
rect 13092 2081 13126 2115
rect 13160 2081 13194 2115
rect 13228 2081 13262 2115
rect 13296 2081 13330 2115
rect 13364 2081 13398 2115
rect 13432 2081 13466 2115
rect 13034 2046 13500 2081
rect 13034 2012 13058 2046
rect 13092 2012 13126 2046
rect 13160 2012 13194 2046
rect 13228 2012 13262 2046
rect 13296 2012 13330 2046
rect 13364 2012 13398 2046
rect 13432 2012 13466 2046
rect 13034 1977 13500 2012
rect 13034 1943 13058 1977
rect 13092 1943 13126 1977
rect 13160 1943 13194 1977
rect 13228 1943 13262 1977
rect 13296 1943 13330 1977
rect 13364 1943 13398 1977
rect 13432 1943 13466 1977
rect 13034 1908 13500 1943
rect 13034 1874 13058 1908
rect 13092 1874 13126 1908
rect 13160 1874 13194 1908
rect 13228 1874 13262 1908
rect 13296 1874 13330 1908
rect 13364 1874 13398 1908
rect 13432 1874 13466 1908
rect 13034 1839 13500 1874
rect 13034 1805 13058 1839
rect 13092 1805 13126 1839
rect 13160 1805 13194 1839
rect 13228 1805 13262 1839
rect 13296 1805 13330 1839
rect 13364 1805 13398 1839
rect 13432 1805 13466 1839
rect 13034 1770 13500 1805
rect 13034 1736 13058 1770
rect 13092 1736 13126 1770
rect 13160 1736 13194 1770
rect 13228 1736 13262 1770
rect 13296 1736 13330 1770
rect 13364 1736 13398 1770
rect 13432 1736 13466 1770
rect 13034 1701 13500 1736
rect 13034 1667 13058 1701
rect 13092 1667 13126 1701
rect 13160 1667 13194 1701
rect 13228 1667 13262 1701
rect 13296 1667 13330 1701
rect 13364 1667 13398 1701
rect 13432 1667 13466 1701
rect 13034 1632 13500 1667
rect 13034 1598 13058 1632
rect 13092 1598 13126 1632
rect 13160 1598 13194 1632
rect 13228 1598 13262 1632
rect 13296 1598 13330 1632
rect 13364 1598 13398 1632
rect 13432 1598 13466 1632
rect 13034 1563 13500 1598
rect 13034 1529 13058 1563
rect 13092 1529 13126 1563
rect 13160 1529 13194 1563
rect 13228 1529 13262 1563
rect 13296 1529 13330 1563
rect 13364 1529 13398 1563
rect 13432 1529 13466 1563
rect 13034 1494 13500 1529
rect 13034 1426 13058 1494
rect 13231 1460 13262 1494
rect 10619 1316 10653 1426
rect 10691 1392 10722 1426
rect 10764 1392 10791 1426
rect 10837 1392 10860 1426
rect 10910 1392 10929 1426
rect 10983 1392 10998 1426
rect 11056 1392 11067 1426
rect 11129 1392 11136 1426
rect 11202 1392 11205 1426
rect 11239 1392 11241 1426
rect 11308 1392 11314 1426
rect 11377 1392 11387 1426
rect 11446 1392 11460 1426
rect 11515 1392 11533 1426
rect 11584 1392 11606 1426
rect 11653 1392 11678 1426
rect 11722 1392 11750 1426
rect 11791 1392 11822 1426
rect 11860 1392 11894 1426
rect 11929 1392 11964 1426
rect 12000 1392 12033 1426
rect 12072 1392 12102 1426
rect 12144 1392 12171 1426
rect 12216 1392 12240 1426
rect 12288 1392 12309 1426
rect 12360 1392 12378 1426
rect 12432 1392 12447 1426
rect 12504 1392 12516 1426
rect 12576 1392 12585 1426
rect 12648 1392 12653 1426
rect 12720 1392 12721 1426
rect 12755 1392 12758 1426
rect 12823 1392 12830 1426
rect 12891 1392 12902 1426
rect 12959 1392 12974 1426
rect 13027 1392 13046 1426
rect 13231 1392 13279 1460
rect 19100 2105 19193 2142
rect 19125 2071 19159 2105
rect 19100 2034 19193 2071
rect 19125 2000 19159 2034
rect 19100 1963 19193 2000
rect 19125 1929 19159 1963
rect 19100 1892 19193 1929
rect 19125 1858 19159 1892
rect 19100 1821 19193 1858
rect 19125 1787 19159 1821
rect 19100 1750 19193 1787
rect 19125 1716 19159 1750
rect 19100 1679 19193 1716
rect 19125 1645 19159 1679
rect 19100 1608 19193 1645
rect 19125 1574 19159 1608
rect 19100 1537 19193 1574
rect 19125 1503 19159 1537
rect 19100 1466 19193 1503
rect 19125 1432 19159 1466
rect 13517 1392 13551 1426
rect 13585 1392 13609 1426
rect 19100 1396 19193 1432
rect 10619 1244 10653 1282
rect 10619 1172 10653 1210
rect 10619 1100 10653 1138
rect 10619 1028 10653 1066
rect 10619 956 10653 994
rect 19125 1362 19159 1396
rect 19100 1326 19193 1362
rect 18994 1292 19091 1301
rect 19125 1292 19159 1326
rect 18994 1262 19193 1292
rect 19028 1228 19066 1262
rect 19100 1256 19193 1262
rect 18994 1222 19091 1228
rect 19125 1222 19159 1256
rect 18994 1189 19193 1222
rect 19028 1155 19066 1189
rect 19100 1186 19193 1189
rect 18994 1152 19091 1155
rect 19125 1152 19159 1186
rect 18994 1116 19193 1152
rect 19028 1082 19066 1116
rect 19125 1082 19159 1116
rect 18994 1046 19193 1082
rect 18994 1043 19091 1046
rect 19028 1009 19066 1043
rect 19125 1012 19159 1046
rect 19100 1009 19193 1012
rect 18994 976 19193 1009
rect 18994 970 19091 976
rect 19028 936 19066 970
rect 19125 942 19159 976
rect 19100 936 19193 942
rect 10619 884 10653 922
rect 19091 918 19193 936
rect 10619 812 10653 850
rect 10619 740 10653 778
rect 10619 668 10653 706
rect 10619 596 10653 634
rect 10619 524 10653 562
rect 10619 452 10653 490
rect 19052 740 19154 764
rect 19086 737 19154 740
rect 19086 706 19114 737
rect 19052 703 19114 706
rect 19148 703 19154 737
rect 19052 667 19154 703
rect 19086 656 19154 667
rect 19086 633 19114 656
rect 19052 622 19114 633
rect 19148 622 19154 656
rect 19052 594 19154 622
rect 19086 575 19154 594
rect 19086 560 19114 575
rect 19052 541 19114 560
rect 19148 541 19154 575
rect 19052 522 19154 541
rect 19086 494 19154 522
rect 19086 488 19114 494
rect 19052 460 19114 488
rect 19148 460 19154 494
rect 19052 450 19154 460
rect 11230 402 11578 436
rect 19086 416 19154 450
rect 19052 413 19154 416
rect 10619 380 10653 394
rect 10619 338 10653 346
rect 19052 379 19114 413
rect 19148 379 19154 413
rect 19052 378 19154 379
rect 19086 344 19154 378
rect 19052 332 19154 344
rect 10653 294 10721 328
rect 10755 294 10790 328
rect 10824 294 10859 328
rect 10893 294 10928 328
rect 10962 294 10997 328
rect 11031 294 11066 328
rect 11100 294 11135 328
rect 11169 294 11204 328
rect 11238 294 11273 328
rect 11307 294 11342 328
rect 11376 294 11411 328
rect 11445 294 11480 328
rect 11514 294 11549 328
rect 11583 294 11618 328
rect 11652 294 11687 328
rect 11721 294 11756 328
rect 11790 294 11825 328
rect 11859 294 11894 328
rect 11928 294 11963 328
rect 11997 294 12032 328
rect 12066 294 12101 328
rect 12135 294 12170 328
rect 12204 294 12239 328
rect 12273 294 12308 328
rect 12342 294 12377 328
rect 12411 294 12446 328
rect 12480 294 12515 328
rect 12549 294 12584 328
rect 12618 294 12653 328
rect 12687 294 12722 328
rect 12756 294 12791 328
rect 12825 294 12860 328
rect 12894 294 12929 328
rect 12963 294 12998 328
rect 13032 294 13067 328
rect 10653 274 13067 294
rect 10619 260 13067 274
rect 10619 248 10721 260
rect 10653 226 10721 248
rect 10755 226 10790 260
rect 10824 226 10859 260
rect 10893 226 10928 260
rect 10962 226 10997 260
rect 11031 226 11066 260
rect 11100 226 11135 260
rect 11169 226 11204 260
rect 11238 226 11273 260
rect 11307 226 11342 260
rect 11376 226 11411 260
rect 11445 226 11480 260
rect 11514 226 11549 260
rect 11583 226 11618 260
rect 11652 226 11687 260
rect 11721 226 11756 260
rect 11790 226 11825 260
rect 11859 226 11894 260
rect 11928 226 11963 260
rect 11997 226 12032 260
rect 12066 226 12101 260
rect 12135 226 12170 260
rect 12204 226 12239 260
rect 12273 226 12308 260
rect 12342 226 12377 260
rect 12411 226 12446 260
rect 12480 226 12515 260
rect 12549 226 12584 260
rect 12618 226 12653 260
rect 12687 226 12722 260
rect 12756 226 12791 260
rect 12825 226 12860 260
rect 12894 226 12929 260
rect 12963 226 12998 260
rect 13032 226 13067 260
rect 10653 201 13067 226
rect 10619 192 13067 201
rect 10619 162 10721 192
rect 10653 158 10721 162
rect 10755 158 10790 192
rect 10824 158 10859 192
rect 10893 158 10928 192
rect 10962 158 10997 192
rect 11031 158 11066 192
rect 11100 158 11135 192
rect 11169 158 11204 192
rect 11238 158 11273 192
rect 11307 158 11342 192
rect 11376 158 11411 192
rect 11445 158 11480 192
rect 11514 158 11549 192
rect 11583 158 11618 192
rect 11652 158 11687 192
rect 11721 158 11756 192
rect 11790 158 11825 192
rect 11859 158 11894 192
rect 11928 158 11963 192
rect 11997 158 12032 192
rect 12066 158 12101 192
rect 12135 158 12170 192
rect 12204 158 12239 192
rect 12273 158 12308 192
rect 12342 158 12377 192
rect 12411 158 12446 192
rect 12480 158 12515 192
rect 12549 158 12584 192
rect 12618 158 12653 192
rect 12687 158 12722 192
rect 12756 158 12791 192
rect 12825 158 12860 192
rect 12894 158 12929 192
rect 12963 158 12998 192
rect 13032 158 13067 192
rect 10653 124 13067 158
rect 15073 294 15097 328
rect 19052 306 19114 332
rect 15073 260 15171 294
rect 15205 260 15240 294
rect 15274 260 15309 294
rect 15343 260 15378 294
rect 15412 260 15447 294
rect 15481 260 15516 294
rect 15550 260 15585 294
rect 15619 260 15654 294
rect 15688 260 15723 294
rect 15757 260 15792 294
rect 15826 260 15861 294
rect 15895 260 15930 294
rect 15964 260 15999 294
rect 16033 260 16068 294
rect 16102 260 16137 294
rect 16171 260 16206 294
rect 16240 260 16275 294
rect 16309 260 16344 294
rect 16378 260 16413 294
rect 16447 260 16482 294
rect 16516 260 16551 294
rect 16585 260 16620 294
rect 16654 260 16689 294
rect 16723 260 16758 294
rect 16792 260 16827 294
rect 16861 260 16896 294
rect 16930 260 16965 294
rect 16999 260 17034 294
rect 17068 260 17103 294
rect 17137 260 17172 294
rect 17206 260 17241 294
rect 17275 260 17310 294
rect 17344 260 17379 294
rect 17413 260 17448 294
rect 17482 260 17517 294
rect 17551 260 17586 294
rect 17620 260 17655 294
rect 17689 260 17724 294
rect 17758 260 17793 294
rect 17827 260 17862 294
rect 17896 260 17931 294
rect 17965 260 18000 294
rect 18034 260 18069 294
rect 18103 260 18138 294
rect 18172 260 18208 294
rect 18242 260 18278 294
rect 18312 260 18348 294
rect 18382 260 18418 294
rect 18452 260 18488 294
rect 18522 260 18558 294
rect 18592 260 18628 294
rect 18662 260 18698 294
rect 18732 260 18768 294
rect 18802 260 18838 294
rect 18872 260 18908 294
rect 18942 260 18978 294
rect 19012 272 19052 294
rect 19086 298 19114 306
rect 19148 298 19154 332
rect 19086 272 19154 298
rect 19012 260 19154 272
rect 15073 251 19154 260
rect 15073 234 19114 251
rect 15073 226 19052 234
rect 15073 192 15171 226
rect 15205 192 15240 226
rect 15274 192 15309 226
rect 15343 192 15378 226
rect 15412 192 15447 226
rect 15481 192 15516 226
rect 15550 192 15585 226
rect 15619 192 15654 226
rect 15688 192 15723 226
rect 15757 192 15792 226
rect 15826 192 15861 226
rect 15895 192 15930 226
rect 15964 192 15999 226
rect 16033 192 16068 226
rect 16102 192 16137 226
rect 16171 192 16206 226
rect 16240 192 16275 226
rect 16309 192 16344 226
rect 16378 192 16413 226
rect 16447 192 16482 226
rect 16516 192 16551 226
rect 16585 192 16620 226
rect 16654 192 16689 226
rect 16723 192 16758 226
rect 16792 192 16827 226
rect 16861 192 16896 226
rect 16930 192 16965 226
rect 16999 192 17034 226
rect 17068 192 17103 226
rect 17137 192 17172 226
rect 17206 192 17241 226
rect 17275 192 17310 226
rect 17344 192 17379 226
rect 17413 192 17448 226
rect 17482 192 17517 226
rect 17551 192 17586 226
rect 17620 192 17655 226
rect 17689 192 17724 226
rect 17758 192 17793 226
rect 17827 192 17862 226
rect 17896 192 17931 226
rect 17965 192 18000 226
rect 18034 192 18069 226
rect 18103 192 18138 226
rect 18172 192 18208 226
rect 18242 192 18278 226
rect 18312 192 18348 226
rect 18382 192 18418 226
rect 18452 192 18488 226
rect 18522 192 18558 226
rect 18592 192 18628 226
rect 18662 192 18698 226
rect 18732 192 18768 226
rect 18802 192 18838 226
rect 18872 192 18908 226
rect 18942 192 18978 226
rect 19012 200 19052 226
rect 19086 217 19114 234
rect 19148 217 19154 251
rect 19086 200 19154 217
rect 19012 192 19154 200
rect 15073 124 19154 192
rect 10619 90 10721 124
rect 10763 90 10789 124
rect 10835 90 10857 124
rect 10907 90 10925 124
rect 10979 90 10993 124
rect 11051 90 11061 124
rect 11123 90 11129 124
rect 11195 90 11197 124
rect 11231 90 11233 124
rect 11299 90 11305 124
rect 11367 90 11377 124
rect 11435 90 11449 124
rect 11503 90 11521 124
rect 11571 90 11593 124
rect 11639 90 11665 124
rect 11707 90 11737 124
rect 11775 90 11809 124
rect 11843 90 11877 124
rect 11915 90 11945 124
rect 11987 90 12013 124
rect 12059 90 12081 124
rect 12131 90 12149 124
rect 12203 90 12217 124
rect 12275 90 12285 124
rect 12347 90 12353 124
rect 12419 90 12421 124
rect 12455 90 12457 124
rect 12523 90 12529 124
rect 12591 90 12601 124
rect 12659 90 12673 124
rect 12727 90 12745 124
rect 12795 90 12817 124
rect 12863 90 12889 124
rect 12931 90 12961 124
rect 12999 90 13033 124
rect 15107 90 15134 124
rect 15175 90 15207 124
rect 15243 90 15277 124
rect 15314 90 15345 124
rect 15387 90 15413 124
rect 15460 90 15481 124
rect 15533 90 15549 124
rect 15606 90 15617 124
rect 15679 90 15685 124
rect 15752 90 15753 124
rect 15787 90 15791 124
rect 15855 90 15864 124
rect 15923 90 15937 124
rect 15991 90 16010 124
rect 16059 90 16083 124
rect 16127 90 16156 124
rect 16195 90 16229 124
rect 16263 90 16297 124
rect 16336 90 16365 124
rect 16409 90 16433 124
rect 16482 90 16501 124
rect 16555 90 16569 124
rect 16628 90 16637 124
rect 16701 90 16705 124
rect 16739 90 16740 124
rect 16807 90 16813 124
rect 16875 90 16886 124
rect 16943 90 16959 124
rect 17011 90 17032 124
rect 17079 90 17105 124
rect 17147 90 17178 124
rect 17215 90 17249 124
rect 17285 90 17317 124
rect 17358 90 17385 124
rect 17431 90 17453 124
rect 17504 90 17521 124
rect 17577 90 17589 124
rect 17650 90 17657 124
rect 17723 90 17725 124
rect 17759 90 17762 124
rect 17827 90 17835 124
rect 17895 90 17908 124
rect 17963 90 17981 124
rect 18031 90 18054 124
rect 18099 90 18127 124
rect 18167 90 18200 124
rect 18235 90 18269 124
rect 18307 90 18337 124
rect 18380 90 18405 124
rect 18453 90 18473 124
rect 18526 90 18541 124
rect 18599 90 18609 124
rect 18672 90 18677 124
rect 18779 90 18784 124
rect 18847 90 18857 124
rect 18915 90 18930 124
rect 18983 90 19003 124
rect 19052 90 19076 124
rect 19110 90 19154 124
rect 18872 64 19154 90
<< viali >>
rect 865 6906 896 6908
rect 896 6906 899 6908
rect 938 6906 965 6908
rect 965 6906 972 6908
rect 1011 6906 1034 6908
rect 1034 6906 1045 6908
rect 1084 6906 1103 6908
rect 1103 6906 1118 6908
rect 1157 6906 1172 6908
rect 1172 6906 1191 6908
rect 1230 6906 1241 6908
rect 1241 6906 1264 6908
rect 1303 6906 1310 6908
rect 1310 6906 1337 6908
rect 1376 6906 1379 6908
rect 1379 6906 1410 6908
rect 1449 6906 1482 6908
rect 1482 6906 1483 6908
rect 1522 6906 1551 6908
rect 1551 6906 1556 6908
rect 1595 6906 1620 6908
rect 1620 6906 1629 6908
rect 1668 6906 1689 6908
rect 1689 6906 1702 6908
rect 1741 6906 1758 6908
rect 1758 6906 1775 6908
rect 1814 6906 1827 6908
rect 1827 6906 1848 6908
rect 865 6874 899 6906
rect 938 6874 972 6906
rect 1011 6874 1045 6906
rect 1084 6874 1118 6906
rect 1157 6874 1191 6906
rect 1230 6874 1264 6906
rect 1303 6874 1337 6906
rect 1376 6874 1410 6906
rect 1449 6874 1483 6906
rect 1522 6874 1556 6906
rect 1595 6874 1629 6906
rect 1668 6874 1702 6906
rect 1741 6874 1775 6906
rect 1814 6874 1848 6906
rect 1887 6874 1921 6908
rect 1960 6874 1994 6908
rect 2033 6874 2067 6908
rect 2106 6874 2140 6908
rect 2179 6874 2213 6908
rect 865 6804 899 6836
rect 938 6804 972 6836
rect 1011 6804 1045 6836
rect 1084 6804 1118 6836
rect 1157 6804 1191 6836
rect 1230 6804 1264 6836
rect 1303 6804 1337 6836
rect 1376 6804 1410 6836
rect 1449 6804 1483 6836
rect 1522 6804 1556 6836
rect 1595 6804 1629 6836
rect 1668 6804 1702 6836
rect 1741 6804 1775 6836
rect 1814 6804 1848 6836
rect 865 6802 896 6804
rect 896 6802 899 6804
rect 938 6802 965 6804
rect 965 6802 972 6804
rect 1011 6802 1034 6804
rect 1034 6802 1045 6804
rect 1084 6802 1103 6804
rect 1103 6802 1118 6804
rect 1157 6802 1172 6804
rect 1172 6802 1191 6804
rect 1230 6802 1241 6804
rect 1241 6802 1264 6804
rect 1303 6802 1310 6804
rect 1310 6802 1337 6804
rect 1376 6802 1379 6804
rect 1379 6802 1410 6804
rect 1449 6802 1482 6804
rect 1482 6802 1483 6804
rect 1522 6802 1551 6804
rect 1551 6802 1556 6804
rect 1595 6802 1620 6804
rect 1620 6802 1629 6804
rect 1668 6802 1689 6804
rect 1689 6802 1702 6804
rect 1741 6802 1758 6804
rect 1758 6802 1775 6804
rect 1814 6802 1827 6804
rect 1827 6802 1848 6804
rect 1887 6802 1921 6836
rect 1960 6802 1994 6836
rect 2033 6802 2067 6836
rect 2106 6802 2140 6836
rect 2179 6802 2213 6836
rect 2252 6802 10056 6908
rect 10056 6906 10090 6908
rect 10090 6906 10124 6908
rect 10124 6906 10158 6908
rect 10158 6906 10192 6908
rect 10192 6906 10226 6908
rect 10226 6906 10260 6908
rect 10260 6906 10294 6908
rect 10294 6906 10328 6908
rect 10328 6906 10362 6908
rect 10362 6906 10396 6908
rect 10396 6906 10430 6908
rect 10430 6906 10464 6908
rect 10464 6906 10498 6908
rect 10498 6906 10532 6908
rect 10532 6906 10566 6908
rect 10566 6906 10600 6908
rect 10600 6906 10634 6908
rect 10634 6906 10668 6908
rect 10668 6906 10702 6908
rect 10702 6906 10736 6908
rect 10736 6906 10770 6908
rect 10770 6906 10804 6908
rect 10804 6906 10838 6908
rect 10838 6906 10872 6908
rect 10872 6906 10906 6908
rect 10906 6906 10940 6908
rect 10940 6906 10974 6908
rect 10974 6906 11008 6908
rect 11008 6906 11042 6908
rect 11042 6906 11076 6908
rect 11076 6906 11110 6908
rect 11110 6906 11144 6908
rect 11144 6906 11178 6908
rect 11178 6906 11212 6908
rect 11212 6906 11246 6908
rect 11246 6906 11280 6908
rect 11280 6906 11314 6908
rect 11314 6906 11348 6908
rect 11348 6906 11382 6908
rect 11382 6906 11416 6908
rect 11416 6906 11450 6908
rect 11450 6906 11484 6908
rect 11484 6906 11518 6908
rect 11518 6906 11552 6908
rect 11552 6906 11586 6908
rect 11586 6906 11620 6908
rect 11620 6906 11654 6908
rect 11654 6906 11688 6908
rect 11688 6906 11722 6908
rect 11722 6906 11756 6908
rect 11756 6906 11790 6908
rect 11790 6906 11824 6908
rect 11824 6906 11858 6908
rect 11858 6906 11892 6908
rect 11892 6906 11926 6908
rect 11926 6906 11960 6908
rect 11960 6906 11994 6908
rect 11994 6906 12028 6908
rect 12028 6906 12062 6908
rect 12062 6906 12096 6908
rect 12096 6906 12130 6908
rect 12130 6906 12164 6908
rect 12164 6906 12198 6908
rect 12198 6906 12232 6908
rect 12232 6906 12266 6908
rect 12266 6906 12300 6908
rect 12300 6906 12334 6908
rect 12334 6906 12368 6908
rect 12368 6906 12402 6908
rect 12402 6906 12436 6908
rect 12436 6906 12471 6908
rect 12471 6906 12505 6908
rect 12505 6906 12540 6908
rect 12540 6906 12574 6908
rect 12574 6906 12609 6908
rect 12609 6906 12643 6908
rect 12643 6906 12678 6908
rect 12678 6906 12712 6908
rect 12712 6906 12747 6908
rect 12747 6906 12781 6908
rect 12781 6906 12816 6908
rect 12816 6906 12850 6908
rect 12850 6906 12885 6908
rect 12885 6906 12919 6908
rect 12919 6906 12954 6908
rect 12954 6906 12988 6908
rect 12988 6906 13023 6908
rect 13023 6906 13057 6908
rect 13057 6906 13092 6908
rect 13092 6906 13126 6908
rect 13126 6906 13161 6908
rect 13161 6906 13195 6908
rect 13195 6906 13230 6908
rect 13230 6906 13264 6908
rect 13264 6906 13299 6908
rect 13299 6906 13302 6908
rect 10056 6872 13302 6906
rect 10056 6838 10091 6872
rect 10091 6838 10125 6872
rect 10125 6838 10160 6872
rect 10160 6838 10194 6872
rect 10194 6838 10229 6872
rect 10229 6838 10263 6872
rect 10263 6838 10298 6872
rect 10298 6838 10332 6872
rect 10332 6838 10367 6872
rect 10367 6838 10401 6872
rect 10401 6838 10436 6872
rect 10436 6838 10470 6872
rect 10470 6838 10505 6872
rect 10505 6838 10539 6872
rect 10539 6838 10574 6872
rect 10574 6838 10608 6872
rect 10608 6838 10643 6872
rect 10643 6838 10677 6872
rect 10677 6838 10712 6872
rect 10712 6838 10746 6872
rect 10746 6838 10781 6872
rect 10781 6838 10815 6872
rect 10815 6838 10850 6872
rect 10850 6838 10884 6872
rect 10884 6838 10919 6872
rect 10919 6838 10953 6872
rect 10953 6838 10988 6872
rect 10988 6838 11022 6872
rect 11022 6838 11057 6872
rect 11057 6838 11091 6872
rect 11091 6838 11126 6872
rect 11126 6838 11160 6872
rect 11160 6838 11195 6872
rect 11195 6838 11229 6872
rect 11229 6838 11264 6872
rect 11264 6838 11298 6872
rect 11298 6838 11333 6872
rect 11333 6838 11367 6872
rect 11367 6838 11402 6872
rect 11402 6838 11436 6872
rect 11436 6838 11471 6872
rect 11471 6838 11505 6872
rect 11505 6838 11540 6872
rect 11540 6838 11574 6872
rect 11574 6838 11609 6872
rect 11609 6838 11643 6872
rect 11643 6838 11678 6872
rect 11678 6838 11712 6872
rect 11712 6838 11747 6872
rect 11747 6838 11781 6872
rect 11781 6838 11816 6872
rect 11816 6838 11850 6872
rect 11850 6838 11885 6872
rect 11885 6838 11919 6872
rect 11919 6838 11954 6872
rect 11954 6838 11988 6872
rect 11988 6838 12023 6872
rect 12023 6838 12057 6872
rect 12057 6838 12092 6872
rect 12092 6838 12126 6872
rect 12126 6838 12161 6872
rect 12161 6838 12195 6872
rect 12195 6838 12230 6872
rect 12230 6838 12264 6872
rect 12264 6838 12299 6872
rect 12299 6838 12333 6872
rect 12333 6838 12368 6872
rect 12368 6838 12402 6872
rect 12402 6838 12437 6872
rect 12437 6838 12471 6872
rect 12471 6838 12506 6872
rect 12506 6838 12540 6872
rect 12540 6838 12575 6872
rect 12575 6838 12609 6872
rect 12609 6838 12644 6872
rect 12644 6838 12678 6872
rect 12678 6838 12713 6872
rect 12713 6838 12747 6872
rect 12747 6838 12782 6872
rect 12782 6838 12816 6872
rect 12816 6838 12851 6872
rect 12851 6838 12885 6872
rect 12885 6838 12920 6872
rect 12920 6838 12954 6872
rect 12954 6838 12989 6872
rect 12989 6838 13023 6872
rect 13023 6838 13058 6872
rect 13058 6838 13092 6872
rect 13092 6838 13127 6872
rect 13127 6838 13161 6872
rect 13161 6838 13196 6872
rect 13196 6838 13230 6872
rect 13230 6838 13265 6872
rect 13265 6838 13299 6872
rect 13299 6838 13302 6872
rect 10056 6804 13265 6838
rect 13265 6804 13302 6838
rect 10056 6802 10091 6804
rect 10091 6802 10125 6804
rect 10125 6802 10160 6804
rect 10160 6802 10194 6804
rect 10194 6802 10229 6804
rect 10229 6802 10263 6804
rect 10263 6802 10298 6804
rect 10298 6802 10332 6804
rect 10332 6802 10367 6804
rect 10367 6802 10401 6804
rect 10401 6802 10436 6804
rect 10436 6802 10470 6804
rect 10470 6802 10505 6804
rect 10505 6802 10539 6804
rect 10539 6802 10574 6804
rect 10574 6802 10608 6804
rect 10608 6802 10643 6804
rect 10643 6802 10677 6804
rect 10677 6802 10712 6804
rect 10712 6802 10746 6804
rect 10746 6802 10781 6804
rect 10781 6802 10815 6804
rect 10815 6802 10850 6804
rect 10850 6802 10884 6804
rect 10884 6802 10919 6804
rect 10919 6802 10953 6804
rect 10953 6802 10988 6804
rect 10988 6802 11022 6804
rect 11022 6802 11057 6804
rect 11057 6802 11091 6804
rect 11091 6802 11126 6804
rect 11126 6802 11160 6804
rect 11160 6802 11195 6804
rect 11195 6802 11229 6804
rect 11229 6802 11264 6804
rect 11264 6802 11298 6804
rect 11298 6802 11333 6804
rect 11333 6802 11367 6804
rect 11367 6802 11402 6804
rect 11402 6802 11436 6804
rect 11436 6802 11471 6804
rect 11471 6802 11505 6804
rect 11505 6802 11540 6804
rect 11540 6802 11574 6804
rect 11574 6802 11609 6804
rect 11609 6802 11643 6804
rect 11643 6802 11678 6804
rect 11678 6802 11712 6804
rect 11712 6802 11747 6804
rect 11747 6802 11781 6804
rect 11781 6802 11816 6804
rect 11816 6802 11850 6804
rect 11850 6802 11885 6804
rect 11885 6802 11919 6804
rect 11919 6802 11954 6804
rect 11954 6802 11988 6804
rect 11988 6802 12023 6804
rect 12023 6802 12057 6804
rect 12057 6802 12092 6804
rect 12092 6802 12126 6804
rect 12126 6802 12161 6804
rect 12161 6802 12195 6804
rect 12195 6802 12230 6804
rect 12230 6802 12264 6804
rect 12264 6802 12299 6804
rect 12299 6802 12333 6804
rect 12333 6802 12368 6804
rect 12368 6802 12402 6804
rect 12402 6802 12437 6804
rect 12437 6802 12471 6804
rect 12471 6802 12506 6804
rect 12506 6802 12540 6804
rect 12540 6802 12575 6804
rect 12575 6802 12609 6804
rect 12609 6802 12644 6804
rect 12644 6802 12678 6804
rect 12678 6802 12713 6804
rect 12713 6802 12747 6804
rect 12747 6802 12782 6804
rect 12782 6802 12816 6804
rect 12816 6802 12851 6804
rect 12851 6802 12885 6804
rect 12885 6802 12920 6804
rect 12920 6802 12954 6804
rect 12954 6802 12989 6804
rect 12989 6802 13023 6804
rect 13023 6802 13058 6804
rect 13058 6802 13092 6804
rect 13092 6802 13127 6804
rect 13127 6802 13161 6804
rect 13161 6802 13197 6804
rect 13197 6764 13302 6804
rect 5870 6633 5904 6667
rect 5945 6633 5979 6667
rect 6020 6633 6054 6667
rect 6095 6633 6129 6667
rect 6170 6633 6204 6667
rect 6245 6633 6279 6667
rect 6319 6633 6353 6667
rect 6393 6633 6427 6667
rect 5792 6538 5826 6563
rect 5792 6529 5826 6538
rect 6522 6538 6556 6563
rect 6522 6529 6556 6538
rect 5792 6470 5826 6491
rect 5792 6457 5826 6470
rect 6522 6470 6556 6491
rect 6522 6457 6556 6470
rect 13197 6730 13303 6764
rect 13197 6657 13231 6691
rect 13269 6657 13303 6691
rect 13197 6584 13231 6618
rect 13269 6584 13303 6618
rect 5870 6377 5904 6411
rect 5945 6377 5979 6411
rect 6020 6377 6054 6411
rect 6095 6377 6129 6411
rect 6170 6377 6204 6411
rect 6245 6377 6279 6411
rect 6319 6377 6353 6411
rect 6393 6377 6427 6411
rect 6932 6289 6966 6323
rect 7005 6289 7039 6323
rect 7078 6289 7112 6323
rect 7151 6289 7185 6323
rect 7224 6289 7258 6323
rect 7297 6289 7331 6323
rect 7370 6289 7404 6323
rect 7443 6289 7477 6323
rect 7516 6289 7550 6323
rect 7589 6289 7623 6323
rect 7662 6289 7696 6323
rect 7735 6289 7769 6323
rect 7808 6289 7842 6323
rect 7881 6289 7915 6323
rect 7954 6289 7988 6323
rect 8027 6289 8061 6323
rect 8100 6289 8134 6323
rect 8173 6289 8207 6323
rect 8246 6289 8280 6323
rect 8319 6289 8353 6323
rect 8392 6289 8426 6323
rect 8465 6289 8499 6323
rect 8538 6289 8572 6323
rect 8611 6289 8645 6323
rect 8684 6289 8718 6323
rect 8757 6289 8791 6323
rect 8830 6289 8864 6323
rect 8903 6289 8937 6323
rect 8976 6289 9010 6323
rect 9049 6289 9083 6323
rect 9122 6289 9156 6323
rect 9195 6289 9229 6323
rect 9268 6289 9302 6323
rect 9341 6289 9375 6323
rect 9414 6289 9448 6323
rect 9486 6289 9520 6323
rect 9558 6289 9592 6323
rect 9630 6289 9664 6323
rect 9702 6289 9736 6323
rect 9774 6289 9808 6323
rect 9846 6289 9880 6323
rect 10131 6289 10165 6323
rect 10203 6289 10237 6323
rect 10275 6289 10309 6323
rect 10347 6289 10381 6323
rect 10419 6289 10453 6323
rect 10491 6289 10525 6323
rect 10563 6289 10597 6323
rect 10635 6289 10669 6323
rect 10707 6289 10741 6323
rect 10779 6289 10813 6323
rect 10852 6289 10886 6323
rect 10925 6289 10959 6323
rect 10998 6289 11032 6323
rect 11071 6289 11105 6323
rect 11144 6289 11178 6323
rect 11217 6289 11251 6323
rect 11290 6289 11324 6323
rect 11363 6289 11397 6323
rect 11436 6289 11470 6323
rect 11509 6289 11543 6323
rect 11582 6289 11616 6323
rect 11655 6289 11689 6323
rect 11728 6289 11762 6323
rect 11801 6289 11835 6323
rect 11874 6289 11908 6323
rect 11947 6289 11981 6323
rect 12020 6289 12054 6323
rect 12093 6289 12127 6323
rect 12166 6289 12200 6323
rect 12239 6289 12273 6323
rect 12312 6289 12346 6323
rect 12385 6289 12419 6323
rect 12458 6289 12492 6323
rect 12531 6289 12565 6323
rect 12604 6289 12638 6323
rect 12677 6289 12711 6323
rect 12750 6289 12784 6323
rect 12823 6289 12857 6323
rect 12896 6289 12930 6323
rect 12969 6289 13003 6323
rect 13042 6289 13076 6323
rect 6852 6279 6886 6281
rect 6852 6247 6886 6279
rect 6852 6177 6886 6209
rect 6852 6175 6886 6177
rect 13122 6279 13156 6281
rect 13122 6247 13125 6279
rect 13125 6247 13156 6279
rect 13122 6177 13125 6209
rect 13125 6177 13156 6209
rect 13122 6175 13156 6177
rect 7172 6133 7206 6167
rect 7246 6133 7280 6167
rect 7320 6133 7354 6167
rect 7394 6133 7428 6167
rect 7468 6133 7502 6167
rect 7542 6133 7576 6167
rect 7616 6133 7650 6167
rect 7690 6133 7724 6167
rect 7764 6133 7798 6167
rect 7837 6133 7871 6167
rect 7910 6133 7944 6167
rect 7983 6133 8017 6167
rect 8056 6133 8090 6167
rect 8129 6133 8163 6167
rect 8202 6133 8236 6167
rect 8275 6133 8309 6167
rect 8348 6133 8382 6167
rect 8421 6133 8455 6167
rect 8494 6133 8528 6167
rect 8567 6133 8601 6167
rect 8640 6133 8674 6167
rect 8713 6133 8747 6167
rect 8786 6133 8820 6167
rect 8859 6133 8893 6167
rect 8932 6133 8966 6167
rect 9005 6133 9039 6167
rect 9078 6133 9112 6167
rect 9151 6133 9185 6167
rect 9224 6133 9258 6167
rect 9297 6133 9331 6167
rect 9370 6133 9404 6167
rect 9443 6133 9477 6167
rect 9516 6133 9550 6167
rect 9589 6133 9623 6167
rect 9662 6133 9696 6167
rect 9735 6133 9769 6167
rect 9808 6133 9842 6167
rect 10169 6133 10203 6167
rect 10242 6133 10276 6167
rect 10315 6133 10349 6167
rect 10388 6133 10422 6167
rect 10461 6133 10495 6167
rect 10534 6133 10568 6167
rect 10607 6133 10641 6167
rect 10680 6133 10714 6167
rect 10753 6133 10787 6167
rect 10826 6133 10860 6167
rect 10899 6133 10933 6167
rect 10972 6133 11006 6167
rect 11045 6133 11079 6167
rect 11118 6133 11152 6167
rect 11191 6133 11225 6167
rect 11264 6133 11298 6167
rect 11337 6133 11371 6167
rect 11410 6133 11444 6167
rect 11483 6133 11517 6167
rect 11556 6133 11590 6167
rect 11629 6133 11663 6167
rect 11702 6133 11736 6167
rect 11775 6133 11809 6167
rect 11848 6133 11882 6167
rect 11921 6133 11955 6167
rect 11994 6133 12028 6167
rect 12067 6133 12101 6167
rect 12140 6133 12174 6167
rect 12213 6133 12247 6167
rect 12286 6133 12320 6167
rect 12359 6133 12393 6167
rect 12432 6133 12466 6167
rect 12506 6133 12540 6167
rect 12580 6133 12614 6167
rect 12654 6133 12688 6167
rect 12728 6133 12762 6167
rect 12802 6133 12836 6167
rect 6932 5941 6966 5975
rect 7005 5941 7039 5975
rect 7078 5941 7112 5975
rect 7151 5941 7185 5975
rect 7224 5941 7258 5975
rect 7297 5941 7331 5975
rect 7370 5941 7404 5975
rect 7443 5941 7477 5975
rect 7516 5941 7550 5975
rect 7589 5941 7623 5975
rect 7662 5941 7696 5975
rect 7735 5941 7769 5975
rect 7808 5941 7842 5975
rect 7881 5941 7915 5975
rect 7954 5941 7988 5975
rect 8027 5941 8061 5975
rect 8100 5941 8134 5975
rect 8173 5941 8207 5975
rect 8246 5941 8280 5975
rect 8319 5941 8353 5975
rect 8392 5941 8426 5975
rect 8465 5941 8499 5975
rect 8538 5941 8572 5975
rect 8611 5941 8645 5975
rect 8684 5941 8718 5975
rect 8757 5941 8791 5975
rect 8830 5941 8864 5975
rect 8903 5941 8937 5975
rect 8976 5941 9010 5975
rect 9049 5941 9083 5975
rect 9122 5941 9156 5975
rect 9195 5941 9229 5975
rect 9268 5941 9302 5975
rect 9341 5941 9375 5975
rect 9414 5941 9448 5975
rect 9486 5941 9520 5975
rect 9558 5941 9592 5975
rect 9630 5941 9664 5975
rect 9702 5941 9736 5975
rect 9774 5941 9808 5975
rect 9846 5941 9880 5975
rect 10131 5941 10165 5975
rect 10203 5941 10237 5975
rect 10275 5941 10309 5975
rect 10347 5941 10381 5975
rect 10419 5941 10453 5975
rect 10491 5941 10525 5975
rect 10563 5941 10597 5975
rect 10635 5941 10669 5975
rect 10707 5941 10741 5975
rect 10779 5941 10813 5975
rect 10852 5941 10886 5975
rect 10925 5941 10959 5975
rect 10998 5941 11032 5975
rect 11071 5941 11105 5975
rect 11144 5941 11178 5975
rect 11217 5941 11251 5975
rect 11290 5941 11324 5975
rect 11363 5941 11397 5975
rect 11436 5941 11470 5975
rect 11509 5941 11543 5975
rect 11582 5941 11616 5975
rect 11655 5941 11689 5975
rect 11728 5941 11762 5975
rect 11801 5941 11835 5975
rect 11874 5941 11908 5975
rect 11947 5941 11981 5975
rect 12020 5941 12054 5975
rect 12093 5941 12127 5975
rect 12166 5941 12200 5975
rect 12239 5941 12273 5975
rect 12312 5941 12346 5975
rect 12385 5941 12419 5975
rect 12458 5941 12492 5975
rect 12531 5941 12565 5975
rect 12604 5941 12638 5975
rect 12677 5941 12711 5975
rect 12750 5941 12784 5975
rect 12823 5941 12857 5975
rect 12896 5941 12930 5975
rect 12969 5941 13003 5975
rect 13042 5941 13076 5975
rect 6852 5930 6886 5931
rect 6852 5897 6886 5930
rect 6852 5828 6886 5859
rect 6852 5825 6886 5828
rect 13122 5931 13156 5933
rect 13122 5899 13125 5931
rect 13125 5899 13156 5931
rect 13122 5829 13125 5861
rect 13125 5829 13156 5861
rect 13122 5827 13156 5829
rect 7181 5785 7215 5819
rect 7254 5785 7288 5819
rect 7327 5785 7361 5819
rect 7400 5785 7434 5819
rect 7473 5785 7507 5819
rect 7546 5785 7580 5819
rect 7619 5785 7653 5819
rect 7692 5785 7726 5819
rect 7765 5785 7799 5819
rect 7838 5785 7872 5819
rect 7911 5785 7945 5819
rect 7984 5785 8018 5819
rect 8057 5785 8091 5819
rect 8130 5785 8164 5819
rect 8203 5785 8237 5819
rect 8276 5785 8310 5819
rect 8349 5785 8383 5819
rect 8422 5785 8456 5819
rect 8494 5785 8528 5819
rect 8566 5785 8600 5819
rect 8638 5785 8672 5819
rect 8710 5785 8744 5819
rect 8782 5785 8816 5819
rect 8854 5785 8888 5819
rect 8926 5785 8960 5819
rect 8998 5785 9032 5819
rect 9070 5785 9104 5819
rect 9142 5785 9176 5819
rect 9214 5785 9248 5819
rect 9286 5785 9320 5819
rect 9358 5785 9392 5819
rect 9430 5785 9464 5819
rect 9502 5785 9536 5819
rect 9574 5785 9608 5819
rect 10169 5785 10203 5819
rect 10242 5785 10276 5819
rect 10315 5785 10349 5819
rect 10388 5785 10422 5819
rect 10461 5785 10495 5819
rect 10534 5785 10568 5819
rect 10607 5785 10641 5819
rect 10680 5785 10714 5819
rect 10753 5785 10787 5819
rect 10826 5785 10860 5819
rect 10899 5785 10933 5819
rect 10972 5785 11006 5819
rect 11045 5785 11079 5819
rect 11118 5785 11152 5819
rect 11191 5785 11225 5819
rect 11264 5785 11298 5819
rect 11337 5785 11371 5819
rect 11410 5785 11444 5819
rect 11483 5785 11517 5819
rect 11556 5785 11590 5819
rect 11629 5785 11663 5819
rect 11702 5785 11736 5819
rect 11775 5785 11809 5819
rect 11848 5785 11882 5819
rect 11921 5785 11955 5819
rect 11994 5785 12028 5819
rect 12067 5785 12101 5819
rect 12140 5785 12174 5819
rect 12213 5785 12247 5819
rect 12286 5785 12320 5819
rect 12359 5785 12393 5819
rect 12432 5785 12466 5819
rect 12506 5785 12540 5819
rect 12580 5785 12614 5819
rect 12654 5785 12688 5819
rect 12728 5785 12762 5819
rect 12802 5785 12836 5819
rect 6932 5593 6966 5627
rect 7005 5593 7039 5627
rect 7078 5593 7112 5627
rect 7151 5593 7185 5627
rect 7224 5593 7258 5627
rect 7297 5593 7331 5627
rect 7370 5593 7404 5627
rect 7443 5593 7477 5627
rect 7516 5593 7550 5627
rect 7589 5593 7623 5627
rect 7662 5593 7696 5627
rect 7735 5593 7769 5627
rect 7808 5593 7842 5627
rect 7881 5593 7915 5627
rect 7954 5593 7988 5627
rect 8027 5593 8061 5627
rect 8100 5593 8134 5627
rect 8173 5593 8207 5627
rect 8246 5593 8280 5627
rect 8319 5593 8353 5627
rect 8392 5593 8426 5627
rect 8465 5593 8499 5627
rect 8538 5593 8572 5627
rect 8611 5593 8645 5627
rect 8684 5593 8718 5627
rect 8757 5593 8791 5627
rect 8830 5593 8864 5627
rect 8903 5593 8937 5627
rect 8976 5593 9010 5627
rect 9049 5593 9083 5627
rect 9122 5593 9156 5627
rect 9195 5593 9229 5627
rect 9268 5593 9302 5627
rect 9341 5593 9375 5627
rect 9414 5593 9448 5627
rect 9486 5593 9520 5627
rect 9558 5593 9592 5627
rect 9630 5593 9664 5627
rect 9702 5593 9736 5627
rect 9774 5593 9808 5627
rect 9846 5593 9880 5627
rect 10131 5593 10165 5627
rect 10203 5593 10237 5627
rect 10275 5593 10309 5627
rect 10347 5593 10381 5627
rect 10419 5593 10453 5627
rect 10491 5593 10525 5627
rect 10563 5593 10597 5627
rect 10635 5593 10669 5627
rect 10707 5593 10741 5627
rect 10779 5593 10813 5627
rect 10852 5593 10886 5627
rect 10925 5593 10959 5627
rect 10998 5593 11032 5627
rect 11071 5593 11105 5627
rect 11144 5593 11178 5627
rect 11217 5593 11251 5627
rect 11290 5593 11324 5627
rect 11363 5593 11397 5627
rect 11436 5593 11470 5627
rect 11509 5593 11543 5627
rect 11582 5593 11616 5627
rect 11655 5593 11689 5627
rect 11728 5593 11762 5627
rect 11801 5593 11835 5627
rect 11874 5593 11908 5627
rect 11947 5593 11981 5627
rect 12020 5593 12054 5627
rect 12093 5593 12127 5627
rect 12166 5593 12200 5627
rect 12239 5593 12273 5627
rect 12312 5593 12346 5627
rect 12385 5593 12419 5627
rect 12458 5593 12492 5627
rect 12531 5593 12565 5627
rect 12604 5593 12638 5627
rect 12677 5593 12711 5627
rect 12750 5593 12784 5627
rect 12823 5593 12857 5627
rect 12896 5593 12930 5627
rect 12969 5593 13003 5627
rect 13042 5593 13076 5627
rect 6852 5583 6886 5584
rect 6852 5550 6886 5583
rect 6852 5481 6886 5512
rect 6852 5478 6886 5481
rect 13122 5583 13156 5585
rect 13122 5551 13125 5583
rect 13125 5551 13156 5583
rect 13122 5481 13125 5513
rect 13125 5481 13156 5513
rect 13122 5479 13156 5481
rect 7172 5437 7206 5471
rect 7246 5437 7280 5471
rect 7320 5437 7354 5471
rect 7394 5437 7428 5471
rect 7468 5437 7502 5471
rect 7542 5437 7576 5471
rect 7616 5437 7650 5471
rect 7690 5437 7724 5471
rect 7764 5437 7798 5471
rect 7838 5437 7872 5471
rect 7912 5437 7946 5471
rect 7985 5437 8019 5471
rect 8058 5437 8092 5471
rect 8131 5437 8165 5471
rect 8204 5437 8238 5471
rect 8277 5437 8311 5471
rect 8350 5437 8384 5471
rect 8423 5437 8457 5471
rect 8496 5437 8530 5471
rect 8569 5437 8603 5471
rect 8642 5437 8676 5471
rect 8715 5437 8749 5471
rect 8788 5437 8822 5471
rect 8861 5437 8895 5471
rect 8934 5437 8968 5471
rect 9007 5437 9041 5471
rect 9080 5437 9114 5471
rect 9153 5437 9187 5471
rect 9226 5437 9260 5471
rect 9299 5437 9333 5471
rect 9372 5437 9406 5471
rect 9445 5437 9479 5471
rect 9518 5437 9552 5471
rect 9591 5437 9625 5471
rect 9664 5437 9698 5471
rect 9737 5437 9771 5471
rect 9810 5437 9844 5471
rect 10169 5437 10203 5471
rect 10242 5437 10276 5471
rect 10315 5437 10349 5471
rect 10388 5437 10422 5471
rect 10461 5437 10495 5471
rect 10534 5437 10568 5471
rect 10607 5437 10641 5471
rect 10680 5437 10714 5471
rect 10753 5437 10787 5471
rect 10826 5437 10860 5471
rect 10899 5437 10933 5471
rect 10972 5437 11006 5471
rect 11045 5437 11079 5471
rect 11118 5437 11152 5471
rect 11191 5437 11225 5471
rect 11264 5437 11298 5471
rect 11337 5437 11371 5471
rect 11410 5437 11444 5471
rect 11483 5437 11517 5471
rect 11556 5437 11590 5471
rect 11629 5437 11663 5471
rect 11702 5437 11736 5471
rect 11775 5437 11809 5471
rect 11848 5437 11882 5471
rect 11921 5437 11955 5471
rect 11994 5437 12028 5471
rect 12067 5437 12101 5471
rect 12140 5437 12174 5471
rect 12213 5437 12247 5471
rect 12286 5437 12320 5471
rect 12359 5437 12393 5471
rect 12432 5437 12466 5471
rect 12506 5437 12540 5471
rect 12580 5437 12614 5471
rect 12654 5437 12688 5471
rect 12728 5437 12762 5471
rect 12802 5437 12836 5471
rect 6932 5245 6966 5279
rect 7005 5245 7039 5279
rect 7078 5245 7112 5279
rect 7151 5245 7185 5279
rect 7224 5245 7258 5279
rect 7297 5245 7331 5279
rect 7370 5245 7404 5279
rect 7443 5245 7477 5279
rect 7516 5245 7550 5279
rect 7589 5245 7623 5279
rect 7662 5245 7696 5279
rect 7735 5245 7769 5279
rect 7808 5245 7842 5279
rect 7881 5245 7915 5279
rect 7954 5245 7988 5279
rect 8027 5245 8061 5279
rect 8100 5245 8134 5279
rect 8173 5245 8207 5279
rect 8246 5245 8280 5279
rect 8319 5245 8353 5279
rect 8392 5245 8426 5279
rect 8465 5245 8499 5279
rect 8538 5245 8572 5279
rect 8611 5245 8645 5279
rect 8684 5245 8718 5279
rect 8757 5245 8791 5279
rect 8830 5245 8864 5279
rect 8903 5245 8937 5279
rect 8976 5245 9010 5279
rect 9049 5245 9083 5279
rect 9122 5245 9156 5279
rect 9195 5245 9229 5279
rect 9268 5245 9302 5279
rect 9341 5245 9375 5279
rect 9414 5245 9448 5279
rect 9486 5245 9520 5279
rect 9558 5245 9592 5279
rect 9630 5245 9664 5279
rect 9702 5245 9736 5279
rect 9774 5245 9808 5279
rect 9846 5245 9880 5279
rect 10131 5245 10165 5279
rect 10203 5245 10237 5279
rect 10275 5245 10309 5279
rect 10347 5245 10381 5279
rect 10419 5245 10453 5279
rect 10491 5245 10525 5279
rect 10563 5245 10597 5279
rect 10635 5245 10669 5279
rect 10707 5245 10741 5279
rect 10779 5245 10813 5279
rect 10852 5245 10886 5279
rect 10925 5245 10959 5279
rect 10998 5245 11032 5279
rect 11071 5245 11105 5279
rect 11144 5245 11178 5279
rect 11217 5245 11251 5279
rect 11290 5245 11324 5279
rect 11363 5245 11397 5279
rect 11436 5245 11470 5279
rect 11509 5245 11543 5279
rect 11582 5245 11616 5279
rect 11655 5245 11689 5279
rect 11728 5245 11762 5279
rect 11801 5245 11835 5279
rect 11874 5245 11908 5279
rect 11947 5245 11981 5279
rect 12020 5245 12054 5279
rect 12093 5245 12127 5279
rect 12166 5245 12200 5279
rect 12239 5245 12273 5279
rect 12312 5245 12346 5279
rect 12385 5245 12419 5279
rect 12458 5245 12492 5279
rect 12531 5245 12565 5279
rect 12604 5245 12638 5279
rect 12677 5245 12711 5279
rect 12750 5245 12784 5279
rect 12823 5245 12857 5279
rect 12896 5245 12930 5279
rect 12969 5245 13003 5279
rect 13042 5245 13076 5279
rect 6852 5235 6886 5244
rect 6852 5210 6886 5235
rect 6852 5167 6886 5172
rect 6852 5138 6886 5167
rect 13122 5235 13156 5252
rect 13122 5218 13125 5235
rect 13125 5218 13156 5235
rect 13122 5167 13156 5180
rect 13122 5146 13125 5167
rect 13125 5146 13156 5167
rect 6932 5089 6966 5123
rect 7006 5089 7040 5123
rect 7080 5089 7114 5123
rect 7154 5089 7188 5123
rect 7228 5089 7262 5123
rect 7302 5089 7336 5123
rect 7376 5089 7410 5123
rect 7450 5089 7484 5123
rect 7524 5089 7558 5123
rect 7597 5089 7631 5123
rect 7670 5089 7704 5123
rect 7743 5089 7777 5123
rect 7816 5089 7850 5123
rect 7889 5089 7923 5123
rect 7962 5089 7996 5123
rect 8035 5089 8069 5123
rect 8108 5089 8142 5123
rect 8181 5089 8215 5123
rect 8254 5089 8288 5123
rect 8327 5089 8361 5123
rect 8400 5089 8434 5123
rect 8473 5089 8507 5123
rect 8546 5089 8580 5123
rect 8619 5089 8653 5123
rect 8692 5089 8726 5123
rect 8765 5089 8799 5123
rect 8838 5089 8872 5123
rect 8911 5089 8945 5123
rect 8984 5089 9018 5123
rect 9057 5089 9091 5123
rect 9130 5089 9164 5123
rect 9203 5089 9237 5123
rect 9276 5089 9310 5123
rect 9349 5089 9383 5123
rect 9422 5089 9456 5123
rect 9495 5089 9529 5123
rect 9568 5089 9602 5123
rect 9641 5089 9675 5123
rect 9714 5089 9748 5123
rect 9787 5089 9821 5123
rect 10196 5089 10230 5123
rect 10268 5089 10302 5123
rect 10341 5089 10375 5123
rect 10414 5089 10448 5123
rect 10487 5089 10521 5123
rect 10560 5089 10594 5123
rect 10633 5089 10667 5123
rect 10706 5089 10740 5123
rect 10779 5089 10813 5123
rect 10852 5089 10886 5123
rect 10925 5089 10959 5123
rect 10998 5089 11032 5123
rect 11071 5089 11105 5123
rect 11144 5089 11178 5123
rect 11217 5089 11251 5123
rect 11290 5089 11324 5123
rect 11363 5089 11397 5123
rect 11436 5089 11470 5123
rect 11509 5089 11543 5123
rect 11582 5089 11616 5123
rect 11655 5089 11689 5123
rect 11728 5089 11762 5123
rect 11801 5089 11835 5123
rect 11874 5089 11908 5123
rect 11947 5089 11981 5123
rect 12020 5089 12054 5123
rect 12093 5089 12127 5123
rect 12166 5089 12200 5123
rect 12239 5089 12273 5123
rect 12312 5089 12346 5123
rect 12385 5089 12419 5123
rect 12458 5089 12492 5123
rect 12531 5089 12565 5123
rect 12604 5089 12638 5123
rect 12677 5089 12711 5123
rect 12750 5089 12784 5123
rect 12823 5089 12857 5123
rect 12896 5089 12930 5123
rect 12969 5089 13003 5123
rect 13042 5089 13076 5123
rect 13197 5143 13303 6545
rect 3410 4729 3443 4731
rect 3443 4729 3444 4731
rect 3483 4729 3512 4731
rect 3512 4729 3517 4731
rect 3556 4729 3581 4731
rect 3581 4729 3590 4731
rect 3629 4729 3650 4731
rect 3650 4729 3663 4731
rect 3702 4729 3719 4731
rect 3719 4729 3736 4731
rect 3775 4729 3788 4731
rect 3788 4729 3809 4731
rect 3848 4729 3857 4731
rect 3857 4729 3882 4731
rect 3921 4729 3926 4731
rect 3926 4729 3955 4731
rect 3994 4729 3995 4731
rect 3995 4729 4028 4731
rect 4067 4729 4098 4731
rect 4098 4729 4101 4731
rect 4140 4729 4167 4731
rect 4167 4729 4174 4731
rect 4213 4729 4236 4731
rect 4236 4729 4247 4731
rect 4286 4729 4305 4731
rect 4305 4729 4320 4731
rect 4359 4729 4374 4731
rect 4374 4729 4393 4731
rect 4432 4729 4443 4731
rect 4443 4729 4466 4731
rect 4505 4729 4512 4731
rect 4512 4729 4539 4731
rect 4578 4729 4581 4731
rect 4581 4729 4612 4731
rect 3410 4697 3444 4729
rect 3483 4697 3517 4729
rect 3556 4697 3590 4729
rect 3629 4697 3663 4729
rect 3702 4697 3736 4729
rect 3775 4697 3809 4729
rect 3848 4697 3882 4729
rect 3921 4697 3955 4729
rect 3994 4697 4028 4729
rect 4067 4697 4101 4729
rect 4140 4697 4174 4729
rect 4213 4697 4247 4729
rect 4286 4697 4320 4729
rect 4359 4697 4393 4729
rect 4432 4697 4466 4729
rect 4505 4697 4539 4729
rect 4578 4697 4612 4729
rect 4651 4697 4685 4731
rect 4724 4729 4754 4731
rect 4754 4729 4758 4731
rect 4797 4729 4823 4731
rect 4823 4729 4831 4731
rect 4870 4729 4892 4731
rect 4892 4729 4904 4731
rect 4943 4729 4961 4731
rect 4961 4729 4977 4731
rect 5016 4729 5030 4731
rect 5030 4729 5050 4731
rect 5089 4729 5099 4731
rect 5099 4729 5123 4731
rect 5162 4729 5168 4731
rect 5168 4729 5196 4731
rect 5235 4729 5237 4731
rect 5237 4729 5269 4731
rect 5307 4729 5340 4731
rect 5340 4729 5341 4731
rect 5379 4729 5409 4731
rect 5409 4729 5413 4731
rect 5451 4729 5478 4731
rect 5478 4729 5485 4731
rect 5523 4729 5547 4731
rect 5547 4729 5557 4731
rect 5595 4729 5616 4731
rect 5616 4729 5629 4731
rect 5667 4729 5685 4731
rect 5685 4729 5701 4731
rect 5739 4729 5754 4731
rect 5754 4729 5773 4731
rect 5811 4729 5823 4731
rect 5823 4729 5845 4731
rect 5883 4729 5892 4731
rect 5892 4729 5917 4731
rect 5955 4729 5961 4731
rect 5961 4729 5989 4731
rect 6027 4729 6030 4731
rect 6030 4729 6061 4731
rect 4724 4697 4758 4729
rect 4797 4697 4831 4729
rect 4870 4697 4904 4729
rect 4943 4697 4977 4729
rect 5016 4697 5050 4729
rect 5089 4697 5123 4729
rect 5162 4697 5196 4729
rect 5235 4697 5269 4729
rect 5307 4697 5341 4729
rect 5379 4697 5413 4729
rect 5451 4697 5485 4729
rect 5523 4697 5557 4729
rect 5595 4697 5629 4729
rect 5667 4697 5701 4729
rect 5739 4697 5773 4729
rect 5811 4697 5845 4729
rect 5883 4697 5917 4729
rect 5955 4697 5989 4729
rect 6027 4697 6061 4729
rect 6099 4697 6133 4731
rect 6171 4729 6203 4731
rect 6203 4729 6205 4731
rect 6243 4729 6272 4731
rect 6272 4729 6277 4731
rect 6315 4729 6341 4731
rect 6341 4729 6349 4731
rect 6387 4729 6410 4731
rect 6410 4729 6421 4731
rect 6459 4729 6479 4731
rect 6479 4729 6493 4731
rect 6531 4729 6548 4731
rect 6548 4729 6565 4731
rect 6603 4729 6617 4731
rect 6617 4729 6637 4731
rect 6675 4729 6686 4731
rect 6686 4729 6709 4731
rect 6747 4729 6755 4731
rect 6755 4729 6781 4731
rect 6819 4729 6824 4731
rect 6824 4729 6853 4731
rect 6891 4729 6893 4731
rect 6893 4729 6925 4731
rect 6171 4697 6205 4729
rect 6243 4697 6277 4729
rect 6315 4697 6349 4729
rect 6387 4697 6421 4729
rect 6459 4697 6493 4729
rect 6531 4697 6565 4729
rect 6603 4697 6637 4729
rect 6675 4697 6709 4729
rect 6747 4697 6781 4729
rect 6819 4697 6853 4729
rect 6891 4697 6925 4729
rect 6963 4697 6997 4731
rect 7035 4697 7069 4731
rect 7107 4697 7141 4731
rect 7179 4697 7213 4731
rect 7251 4697 7285 4731
rect 7323 4697 7357 4731
rect 7395 4697 7429 4731
rect 7467 4697 7501 4731
rect 7539 4697 7573 4731
rect 7611 4697 7645 4731
rect 7683 4697 7717 4731
rect 7755 4697 7789 4731
rect 7827 4697 7861 4731
rect 7899 4697 7933 4731
rect 7971 4697 8005 4731
rect 3444 4627 3478 4659
rect 3517 4627 3551 4659
rect 3590 4627 3624 4659
rect 3663 4627 3697 4659
rect 3736 4627 3770 4659
rect 3809 4627 3843 4659
rect 3882 4627 3916 4659
rect 3955 4627 3989 4659
rect 4028 4627 4062 4659
rect 4101 4627 4135 4659
rect 4174 4627 4208 4659
rect 4247 4627 4281 4659
rect 4320 4627 4354 4659
rect 4393 4627 4427 4659
rect 4466 4627 4500 4659
rect 4539 4627 4573 4659
rect 4612 4627 4646 4659
rect 3444 4625 3476 4627
rect 3476 4625 3478 4627
rect 3517 4625 3545 4627
rect 3545 4625 3551 4627
rect 3590 4625 3614 4627
rect 3614 4625 3624 4627
rect 3663 4625 3683 4627
rect 3683 4625 3697 4627
rect 3736 4625 3752 4627
rect 3752 4625 3770 4627
rect 3809 4625 3821 4627
rect 3821 4625 3843 4627
rect 3882 4625 3890 4627
rect 3890 4625 3916 4627
rect 3955 4625 3959 4627
rect 3959 4625 3989 4627
rect 3372 4587 3406 4613
rect 4028 4625 4062 4627
rect 4101 4625 4131 4627
rect 4131 4625 4135 4627
rect 4174 4625 4200 4627
rect 4200 4625 4208 4627
rect 4247 4625 4269 4627
rect 4269 4625 4281 4627
rect 4320 4625 4338 4627
rect 4338 4625 4354 4627
rect 4393 4625 4407 4627
rect 4407 4625 4427 4627
rect 4466 4625 4476 4627
rect 4476 4625 4500 4627
rect 4539 4625 4545 4627
rect 4545 4625 4573 4627
rect 4612 4625 4614 4627
rect 4614 4625 4646 4627
rect 4685 4625 4718 4659
rect 4718 4625 4719 4659
rect 4758 4625 4792 4659
rect 4831 4625 4865 4659
rect 4904 4625 4938 4659
rect 4977 4625 5011 4659
rect 5050 4625 5084 4659
rect 5123 4625 5157 4659
rect 5196 4625 5230 4659
rect 5269 4625 5303 4659
rect 5342 4625 5376 4659
rect 5415 4625 5449 4659
rect 5488 4625 5522 4659
rect 5561 4625 5595 4659
rect 5634 4625 5668 4659
rect 5707 4625 5741 4659
rect 5780 4625 5814 4659
rect 5853 4625 5887 4659
rect 5926 4625 5960 4659
rect 5999 4625 6033 4659
rect 6072 4625 6106 4659
rect 6145 4625 6179 4659
rect 6218 4625 6252 4659
rect 6291 4625 6325 4659
rect 6364 4625 6398 4659
rect 6437 4625 6471 4659
rect 6510 4625 6544 4659
rect 6583 4625 6617 4659
rect 6656 4625 6690 4659
rect 6729 4625 6763 4659
rect 6802 4625 6836 4659
rect 6875 4625 6909 4659
rect 6948 4625 6982 4659
rect 7021 4625 7055 4659
rect 7094 4625 7128 4659
rect 7167 4625 7201 4659
rect 7240 4625 7274 4659
rect 7313 4625 7347 4659
rect 7386 4625 7420 4659
rect 7459 4625 7493 4659
rect 7532 4625 7566 4659
rect 7605 4625 7639 4659
rect 7678 4625 7712 4659
rect 7751 4625 7785 4659
rect 7824 4625 7858 4659
rect 7897 4625 7931 4659
rect 7970 4625 8004 4659
rect 8043 4625 10056 4731
rect 10056 4729 10092 4731
rect 10092 4729 10126 4731
rect 10126 4729 10161 4731
rect 10161 4729 10195 4731
rect 10195 4729 10230 4731
rect 10230 4729 10264 4731
rect 10264 4729 10299 4731
rect 10299 4729 10333 4731
rect 10333 4729 10368 4731
rect 10368 4729 10402 4731
rect 10402 4729 10437 4731
rect 10437 4729 10471 4731
rect 10471 4729 10506 4731
rect 10506 4729 10540 4731
rect 10540 4729 10575 4731
rect 10575 4729 10609 4731
rect 10609 4729 10644 4731
rect 10644 4729 10678 4731
rect 10678 4729 10713 4731
rect 10713 4729 10747 4731
rect 10747 4729 10782 4731
rect 10782 4729 10816 4731
rect 10816 4729 10851 4731
rect 10851 4729 10885 4731
rect 10885 4729 10920 4731
rect 10920 4729 10954 4731
rect 10954 4729 10989 4731
rect 10989 4729 11023 4731
rect 11023 4729 11058 4731
rect 11058 4729 11092 4731
rect 11092 4729 11127 4731
rect 11127 4729 11161 4731
rect 11161 4729 11196 4731
rect 11196 4729 11230 4731
rect 11230 4729 11265 4731
rect 11265 4729 11299 4731
rect 11299 4729 11334 4731
rect 11334 4729 11368 4731
rect 11368 4729 11403 4731
rect 11403 4729 11437 4731
rect 11437 4729 11472 4731
rect 11472 4729 11506 4731
rect 11506 4729 11541 4731
rect 11541 4729 11575 4731
rect 11575 4729 11610 4731
rect 11610 4729 11644 4731
rect 11644 4729 11679 4731
rect 11679 4729 11713 4731
rect 11713 4729 11748 4731
rect 11748 4729 11782 4731
rect 11782 4729 11817 4731
rect 11817 4729 11851 4731
rect 11851 4729 11886 4731
rect 11886 4729 11920 4731
rect 11920 4729 11955 4731
rect 11955 4729 11989 4731
rect 11989 4729 12024 4731
rect 12024 4729 12058 4731
rect 12058 4729 12093 4731
rect 12093 4729 12127 4731
rect 12127 4729 12162 4731
rect 12162 4729 12196 4731
rect 12196 4729 12231 4731
rect 12231 4729 12265 4731
rect 12265 4729 12300 4731
rect 12300 4729 12334 4731
rect 12334 4729 12369 4731
rect 12369 4729 12403 4731
rect 12403 4729 12438 4731
rect 12438 4729 12472 4731
rect 12472 4729 12507 4731
rect 12507 4729 12541 4731
rect 12541 4729 12576 4731
rect 12576 4729 12610 4731
rect 12610 4729 12645 4731
rect 12645 4729 12679 4731
rect 12679 4729 12714 4731
rect 12714 4729 12748 4731
rect 12748 4729 12783 4731
rect 12783 4729 12817 4731
rect 12817 4729 12852 4731
rect 12852 4729 12886 4731
rect 12886 4729 12921 4731
rect 12921 4729 12955 4731
rect 12955 4729 12990 4731
rect 12990 4729 13024 4731
rect 13024 4729 13059 4731
rect 13059 4729 13093 4731
rect 13093 4729 13128 4731
rect 13128 4729 13162 4731
rect 13162 4729 13197 4731
rect 13197 4729 13231 4731
rect 13231 4730 13265 4731
rect 13265 4730 13333 4731
rect 13231 4729 13333 4730
rect 10056 4695 13333 4729
rect 10056 4661 10091 4695
rect 10091 4661 10125 4695
rect 10125 4661 10160 4695
rect 10160 4661 10194 4695
rect 10194 4661 10229 4695
rect 10229 4661 10263 4695
rect 10263 4661 10298 4695
rect 10298 4661 10332 4695
rect 10332 4661 10367 4695
rect 10367 4661 10401 4695
rect 10401 4661 10436 4695
rect 10436 4661 10470 4695
rect 10470 4661 10505 4695
rect 10505 4661 10539 4695
rect 10539 4661 10574 4695
rect 10574 4661 10608 4695
rect 10608 4661 10643 4695
rect 10643 4661 10677 4695
rect 10677 4661 10712 4695
rect 10712 4661 10746 4695
rect 10746 4661 10781 4695
rect 10781 4661 10815 4695
rect 10815 4661 10850 4695
rect 10850 4661 10884 4695
rect 10884 4661 10919 4695
rect 10919 4661 10953 4695
rect 10953 4661 10988 4695
rect 10988 4661 11022 4695
rect 11022 4661 11057 4695
rect 11057 4661 11091 4695
rect 11091 4661 11126 4695
rect 11126 4661 11160 4695
rect 11160 4661 11195 4695
rect 11195 4661 11229 4695
rect 11229 4661 11264 4695
rect 11264 4661 11298 4695
rect 11298 4661 11333 4695
rect 11333 4661 11367 4695
rect 11367 4661 11402 4695
rect 11402 4661 11436 4695
rect 11436 4661 11471 4695
rect 11471 4661 11505 4695
rect 11505 4661 11540 4695
rect 11540 4661 11574 4695
rect 11574 4661 11609 4695
rect 11609 4661 11643 4695
rect 11643 4661 11678 4695
rect 11678 4661 11712 4695
rect 11712 4661 11747 4695
rect 11747 4661 11781 4695
rect 11781 4661 11816 4695
rect 11816 4661 11850 4695
rect 11850 4661 11885 4695
rect 11885 4661 11919 4695
rect 11919 4661 11954 4695
rect 11954 4661 11988 4695
rect 11988 4661 12023 4695
rect 12023 4661 12057 4695
rect 12057 4661 12092 4695
rect 12092 4661 12126 4695
rect 12126 4661 12161 4695
rect 12161 4661 12195 4695
rect 12195 4661 12230 4695
rect 12230 4661 12264 4695
rect 12264 4661 12299 4695
rect 12299 4661 12333 4695
rect 12333 4661 12368 4695
rect 12368 4661 12402 4695
rect 12402 4661 12437 4695
rect 12437 4661 12471 4695
rect 12471 4661 12506 4695
rect 12506 4661 12540 4695
rect 12540 4661 12575 4695
rect 12575 4661 12609 4695
rect 12609 4661 12644 4695
rect 12644 4661 12678 4695
rect 12678 4661 12713 4695
rect 12713 4661 12747 4695
rect 12747 4661 12782 4695
rect 12782 4661 12816 4695
rect 12816 4661 12851 4695
rect 12851 4661 12885 4695
rect 12885 4661 12920 4695
rect 12920 4661 12954 4695
rect 12954 4661 12989 4695
rect 12989 4661 13023 4695
rect 13023 4661 13058 4695
rect 13058 4661 13092 4695
rect 13092 4661 13127 4695
rect 13127 4661 13161 4695
rect 13161 4661 13196 4695
rect 13196 4661 13230 4695
rect 13230 4661 13265 4695
rect 13265 4661 13299 4695
rect 13299 4661 13333 4695
rect 10056 4627 13333 4661
rect 10056 4625 10091 4627
rect 10091 4625 10125 4627
rect 10125 4625 10160 4627
rect 10160 4625 10194 4627
rect 10194 4625 10229 4627
rect 10229 4625 10263 4627
rect 10263 4625 10298 4627
rect 10298 4625 10332 4627
rect 10332 4625 10367 4627
rect 10367 4625 10401 4627
rect 10401 4625 10436 4627
rect 10436 4625 10470 4627
rect 10470 4625 10505 4627
rect 10505 4625 10539 4627
rect 10539 4625 10574 4627
rect 10574 4625 10608 4627
rect 10608 4625 10643 4627
rect 10643 4625 10677 4627
rect 10677 4625 10712 4627
rect 10712 4625 10746 4627
rect 10746 4625 10781 4627
rect 10781 4625 10815 4627
rect 10815 4625 10850 4627
rect 10850 4625 10884 4627
rect 10884 4625 10919 4627
rect 10919 4625 10953 4627
rect 10953 4625 10987 4627
rect 10987 4625 11021 4627
rect 11021 4625 11055 4627
rect 11055 4625 11089 4627
rect 11089 4625 11123 4627
rect 11123 4625 11157 4627
rect 11157 4625 11191 4627
rect 11191 4625 11225 4627
rect 11225 4625 11259 4627
rect 11259 4625 11293 4627
rect 11293 4625 11327 4627
rect 11327 4625 11361 4627
rect 11361 4625 11395 4627
rect 11395 4625 11429 4627
rect 11429 4625 11463 4627
rect 11463 4625 11497 4627
rect 11497 4625 11531 4627
rect 11531 4625 11565 4627
rect 11565 4625 11599 4627
rect 11599 4625 11633 4627
rect 11633 4625 11667 4627
rect 11667 4625 11701 4627
rect 11701 4625 11735 4627
rect 11735 4625 11769 4627
rect 11769 4625 11803 4627
rect 11803 4625 11837 4627
rect 11837 4625 11871 4627
rect 11871 4625 11905 4627
rect 11905 4625 11939 4627
rect 11939 4625 11973 4627
rect 11973 4625 12007 4627
rect 12007 4625 12041 4627
rect 12041 4625 12075 4627
rect 12075 4625 12109 4627
rect 12109 4625 12143 4627
rect 12143 4625 12177 4627
rect 12177 4625 12211 4627
rect 12211 4625 12245 4627
rect 12245 4625 12279 4627
rect 12279 4625 12313 4627
rect 12313 4625 12347 4627
rect 12347 4625 12381 4627
rect 12381 4625 12415 4627
rect 12415 4625 12449 4627
rect 12449 4625 12483 4627
rect 12483 4625 12517 4627
rect 12517 4625 12551 4627
rect 12551 4625 12585 4627
rect 12585 4625 12619 4627
rect 12619 4625 12653 4627
rect 12653 4625 12687 4627
rect 12687 4625 12721 4627
rect 12721 4625 12755 4627
rect 12755 4625 12789 4627
rect 12789 4625 12823 4627
rect 12823 4625 12857 4627
rect 12857 4625 12891 4627
rect 12891 4625 12925 4627
rect 12925 4625 12959 4627
rect 12959 4625 12993 4627
rect 12993 4625 13027 4627
rect 13027 4625 13061 4627
rect 13061 4625 13095 4627
rect 13095 4625 13129 4627
rect 13129 4625 13163 4627
rect 13163 4625 13197 4627
rect 13197 4625 13231 4627
rect 13231 4625 13265 4627
rect 13265 4625 13333 4627
rect 3372 4579 3374 4587
rect 3374 4579 3406 4587
rect 3444 4557 3478 4582
rect 3372 4517 3406 4537
rect 3372 4503 3374 4517
rect 3374 4503 3406 4517
rect 3444 4548 3476 4557
rect 3476 4548 3478 4557
rect 3444 4487 3478 4505
rect 3372 4447 3406 4461
rect 3372 4427 3374 4447
rect 3374 4427 3406 4447
rect 3444 4471 3476 4487
rect 3476 4471 3478 4487
rect 3444 4417 3478 4428
rect 3372 4377 3406 4384
rect 3372 4350 3374 4377
rect 3374 4350 3406 4377
rect 3444 4394 3476 4417
rect 3476 4394 3478 4417
rect 3444 4347 3478 4351
rect 3372 4273 3374 4307
rect 3374 4273 3406 4307
rect 3444 4317 3476 4347
rect 3476 4317 3478 4347
rect 3372 4203 3374 4230
rect 3374 4203 3406 4230
rect 3444 4243 3476 4274
rect 3476 4243 3478 4274
rect 3444 4240 3478 4243
rect 3372 4196 3406 4203
rect 3372 4133 3374 4153
rect 3374 4133 3406 4153
rect 3444 4173 3476 4197
rect 3476 4173 3478 4197
rect 3444 4163 3478 4173
rect 3372 4119 3406 4133
rect 3372 4062 3374 4076
rect 3374 4062 3406 4076
rect 3444 4102 3476 4120
rect 3476 4102 3478 4120
rect 3444 4086 3478 4102
rect 16111 4142 16145 4176
rect 16111 4070 16145 4104
rect 16287 4142 16321 4176
rect 16287 4070 16321 4104
rect 16463 4142 16497 4176
rect 16463 4070 16497 4104
rect 16639 4142 16673 4176
rect 16639 4070 16673 4104
rect 16837 4142 16871 4176
rect 16837 4070 16871 4104
rect 3372 4042 3406 4062
rect 3444 4031 3476 4043
rect 3476 4031 3478 4043
rect 3444 4009 3478 4031
rect 3372 3991 3374 3999
rect 3374 3991 3406 3999
rect 3372 3965 3406 3991
rect 3444 3960 3476 3966
rect 3476 3960 3478 3966
rect 3444 3932 3478 3960
rect 35 3920 68 3922
rect 68 3920 69 3922
rect 108 3920 137 3922
rect 137 3920 142 3922
rect 181 3920 206 3922
rect 206 3920 215 3922
rect 254 3920 275 3922
rect 275 3920 288 3922
rect 327 3920 344 3922
rect 344 3920 361 3922
rect 400 3920 413 3922
rect 413 3920 434 3922
rect 473 3920 482 3922
rect 482 3920 507 3922
rect 546 3920 551 3922
rect 551 3920 580 3922
rect 35 3888 69 3920
rect 108 3888 142 3920
rect 181 3888 215 3920
rect 254 3888 288 3920
rect 327 3888 361 3920
rect 400 3888 434 3920
rect 473 3888 507 3920
rect 546 3888 580 3920
rect 619 3888 620 3922
rect 620 3888 653 3922
rect 692 3888 726 3922
rect 765 3888 799 3922
rect 838 3888 872 3922
rect 911 3888 945 3922
rect 984 3888 1018 3922
rect 1057 3888 1091 3922
rect 1130 3888 1164 3922
rect 1203 3888 1237 3922
rect 1276 3888 1310 3922
rect 1349 3888 1383 3922
rect 1422 3888 1456 3922
rect 1495 3888 1529 3922
rect 1568 3888 1602 3922
rect 1641 3888 1675 3922
rect 1714 3888 1748 3922
rect 1787 3888 1821 3922
rect 1860 3888 1894 3922
rect 1932 3888 1966 3922
rect 2004 3888 2038 3922
rect 2076 3888 2110 3922
rect 2148 3888 2182 3922
rect 2220 3888 2254 3922
rect 2292 3888 2326 3922
rect 2364 3888 2398 3922
rect 2436 3888 2470 3922
rect 2508 3888 2542 3922
rect 2580 3888 2614 3922
rect 2652 3888 2686 3922
rect 2724 3888 2758 3922
rect 2796 3888 2830 3922
rect 2868 3888 2902 3922
rect 2940 3888 2974 3922
rect 3012 3888 3046 3922
rect 3084 3888 3118 3922
rect 3156 3888 3190 3922
rect 3228 3888 3262 3922
rect 3300 3888 3334 3922
rect 3372 3888 3374 3922
rect 3374 3888 3406 3922
rect 3444 3854 3478 3888
rect 35 3818 69 3850
rect 109 3818 143 3850
rect 183 3818 217 3850
rect 257 3818 291 3850
rect 331 3818 365 3850
rect 405 3818 439 3850
rect 479 3818 513 3850
rect 553 3818 587 3850
rect 627 3818 661 3850
rect 701 3818 735 3850
rect 775 3818 809 3850
rect 849 3818 883 3850
rect 923 3818 957 3850
rect 996 3818 1030 3850
rect 35 3816 68 3818
rect 68 3816 69 3818
rect 109 3816 137 3818
rect 137 3816 143 3818
rect 183 3816 206 3818
rect 206 3816 217 3818
rect 257 3816 275 3818
rect 275 3816 291 3818
rect 331 3816 344 3818
rect 344 3816 365 3818
rect 405 3816 413 3818
rect 413 3816 439 3818
rect 479 3816 482 3818
rect 482 3816 513 3818
rect 553 3816 585 3818
rect 585 3816 587 3818
rect 627 3816 654 3818
rect 654 3816 661 3818
rect 701 3816 723 3818
rect 723 3816 735 3818
rect 775 3816 792 3818
rect 792 3816 809 3818
rect 849 3816 861 3818
rect 861 3816 883 3818
rect 923 3816 930 3818
rect 930 3816 957 3818
rect 996 3816 999 3818
rect 999 3816 1030 3818
rect 1069 3816 1103 3850
rect 1142 3818 1176 3850
rect 1215 3818 1249 3850
rect 1288 3818 1322 3850
rect 1361 3818 1395 3850
rect 1434 3818 1468 3850
rect 1507 3818 1541 3850
rect 1580 3818 1614 3850
rect 1653 3818 1687 3850
rect 1726 3818 1760 3850
rect 1799 3818 1833 3850
rect 1872 3818 1906 3850
rect 1945 3818 1979 3850
rect 2018 3818 2052 3850
rect 2091 3818 2125 3850
rect 2164 3818 2198 3850
rect 2237 3818 2271 3850
rect 1142 3816 1172 3818
rect 1172 3816 1176 3818
rect 1215 3816 1241 3818
rect 1241 3816 1249 3818
rect 1288 3816 1310 3818
rect 1310 3816 1322 3818
rect 1361 3816 1379 3818
rect 1379 3816 1395 3818
rect 1434 3816 1448 3818
rect 1448 3816 1468 3818
rect 1507 3816 1517 3818
rect 1517 3816 1541 3818
rect 1580 3816 1586 3818
rect 1586 3816 1614 3818
rect 1653 3816 1655 3818
rect 1655 3816 1687 3818
rect 1726 3816 1758 3818
rect 1758 3816 1760 3818
rect 1799 3816 1827 3818
rect 1827 3816 1833 3818
rect 1872 3816 1896 3818
rect 1896 3816 1906 3818
rect 1945 3816 1965 3818
rect 1965 3816 1979 3818
rect 2018 3816 2034 3818
rect 2034 3816 2052 3818
rect 2091 3816 2103 3818
rect 2103 3816 2125 3818
rect 2164 3816 2172 3818
rect 2172 3816 2198 3818
rect 2237 3816 2241 3818
rect 2241 3816 2271 3818
rect 2310 3816 2344 3850
rect 2383 3818 2417 3850
rect 2456 3818 2490 3850
rect 2529 3818 2563 3850
rect 2602 3818 2636 3850
rect 2675 3818 2709 3850
rect 2748 3818 2782 3850
rect 2821 3818 2855 3850
rect 2894 3818 2928 3850
rect 2383 3816 2414 3818
rect 2414 3816 2417 3818
rect 2456 3816 2483 3818
rect 2483 3816 2490 3818
rect 2529 3816 2552 3818
rect 2552 3816 2563 3818
rect 2602 3816 2621 3818
rect 2621 3816 2636 3818
rect 2675 3816 2690 3818
rect 2690 3816 2709 3818
rect 2748 3816 2759 3818
rect 2759 3816 2782 3818
rect 2821 3816 2828 3818
rect 2828 3816 2855 3818
rect 2894 3816 2897 3818
rect 2897 3816 2928 3818
rect 2967 3816 3001 3850
rect 3040 3816 3074 3850
rect 3113 3816 3147 3850
rect 3186 3816 3220 3850
rect 3259 3816 3293 3850
rect 3332 3816 3366 3850
rect 16199 3686 16233 3720
rect 16551 3686 16585 3720
rect 16924 3684 16958 3718
rect 16924 3612 16958 3646
rect 13425 3103 13459 3137
rect 13498 3103 13532 3137
rect 13571 3103 13605 3137
rect 13644 3103 13678 3137
rect 13717 3103 13751 3137
rect 13790 3103 13824 3137
rect 13863 3103 13897 3137
rect 13936 3103 13970 3137
rect 14009 3103 14043 3137
rect 14082 3103 14116 3137
rect 14155 3103 14189 3137
rect 14228 3103 14262 3137
rect 14301 3103 14335 3137
rect 14374 3103 14408 3137
rect 14447 3103 14481 3137
rect 14519 3103 14553 3137
rect 14591 3103 14625 3137
rect 14663 3103 14697 3137
rect 14735 3103 14769 3137
rect 14807 3103 14841 3137
rect 14879 3103 14913 3137
rect 14951 3103 14985 3137
rect 15023 3103 15057 3137
rect 15095 3103 15129 3137
rect 15167 3103 15201 3137
rect 15239 3103 15273 3137
rect 15311 3103 15345 3137
rect 15383 3103 15417 3137
rect 15455 3103 15489 3137
rect 15527 3103 15561 3137
rect 15599 3103 15633 3137
rect 15671 3103 15705 3137
rect 15743 3103 15777 3137
rect 15815 3103 15849 3137
rect 15887 3103 15921 3137
rect 15959 3103 15993 3137
rect 16031 3103 16065 3137
rect 16103 3103 16137 3137
rect 16175 3103 16209 3137
rect 16247 3103 16281 3137
rect 16319 3103 16353 3137
rect 16391 3103 16425 3137
rect 16463 3103 16497 3137
rect 16535 3103 16569 3137
rect 16607 3103 16641 3137
rect 16679 3103 16713 3137
rect 16751 3103 16785 3137
rect 16823 3103 16857 3137
rect 16895 3103 16929 3137
rect 16967 3103 17001 3137
rect 17039 3103 17073 3137
rect 17111 3103 17145 3137
rect 17183 3103 17217 3137
rect 17255 3103 17289 3137
rect 17327 3103 17361 3137
rect 17399 3103 17433 3137
rect 17471 3103 17505 3137
rect 17543 3103 17577 3137
rect 17615 3103 17649 3137
rect 17687 3103 17721 3137
rect 17759 3103 17793 3137
rect 17831 3103 17865 3137
rect 17903 3103 17937 3137
rect 17975 3103 18009 3137
rect 18047 3103 18081 3137
rect 18119 3103 18153 3137
rect 18191 3103 18225 3137
rect 18263 3103 18297 3137
rect 18335 3103 18369 3137
rect 18407 3103 18441 3137
rect 18479 3103 18513 3137
rect 18551 3103 18585 3137
rect 18623 3103 18657 3137
rect 18695 3103 18729 3137
rect 18767 3103 18801 3137
rect 18839 3103 18873 3137
rect 18911 3103 18945 3137
rect 18983 3103 19017 3137
rect 19093 3065 19127 3099
rect 19093 2989 19127 3023
rect 19093 2945 19127 2947
rect 19093 2913 19127 2945
rect 19093 2841 19127 2872
rect 19093 2838 19127 2841
rect 19093 2772 19127 2797
rect 19093 2763 19127 2772
rect 19093 2703 19127 2722
rect 19093 2688 19127 2703
rect 19093 2634 19127 2647
rect 19093 2613 19127 2634
rect 19093 2565 19127 2572
rect 19093 2538 19127 2565
rect 19093 2496 19127 2497
rect 19093 2463 19127 2496
rect 18994 2247 19100 2271
rect 18994 2213 19091 2247
rect 19091 2213 19100 2247
rect 18994 2176 19100 2213
rect 18994 2142 19091 2176
rect 19091 2142 19100 2176
rect 10657 1392 10687 1426
rect 10687 1392 10691 1426
rect 10730 1392 10756 1426
rect 10756 1392 10764 1426
rect 10803 1392 10825 1426
rect 10825 1392 10837 1426
rect 10876 1392 10894 1426
rect 10894 1392 10910 1426
rect 10949 1392 10963 1426
rect 10963 1392 10983 1426
rect 11022 1392 11032 1426
rect 11032 1392 11056 1426
rect 11095 1392 11101 1426
rect 11101 1392 11129 1426
rect 11168 1392 11170 1426
rect 11170 1392 11202 1426
rect 11241 1392 11274 1426
rect 11274 1392 11275 1426
rect 11314 1392 11343 1426
rect 11343 1392 11348 1426
rect 11387 1392 11412 1426
rect 11412 1392 11421 1426
rect 11460 1392 11481 1426
rect 11481 1392 11494 1426
rect 11533 1392 11550 1426
rect 11550 1392 11567 1426
rect 11606 1392 11619 1426
rect 11619 1392 11640 1426
rect 11678 1392 11688 1426
rect 11688 1392 11712 1426
rect 11750 1392 11757 1426
rect 11757 1392 11784 1426
rect 11822 1392 11826 1426
rect 11826 1392 11856 1426
rect 11894 1392 11895 1426
rect 11895 1392 11928 1426
rect 11966 1392 11998 1426
rect 11998 1392 12000 1426
rect 12038 1392 12067 1426
rect 12067 1392 12072 1426
rect 12110 1392 12136 1426
rect 12136 1392 12144 1426
rect 12182 1392 12205 1426
rect 12205 1392 12216 1426
rect 12254 1392 12274 1426
rect 12274 1392 12288 1426
rect 12326 1392 12343 1426
rect 12343 1392 12360 1426
rect 12398 1392 12412 1426
rect 12412 1392 12432 1426
rect 12470 1392 12481 1426
rect 12481 1392 12504 1426
rect 12542 1392 12550 1426
rect 12550 1392 12576 1426
rect 12614 1392 12619 1426
rect 12619 1392 12648 1426
rect 12686 1392 12687 1426
rect 12687 1392 12720 1426
rect 12758 1392 12789 1426
rect 12789 1392 12792 1426
rect 12830 1392 12857 1426
rect 12857 1392 12864 1426
rect 12902 1392 12925 1426
rect 12925 1392 12936 1426
rect 12974 1392 12993 1426
rect 12993 1392 13008 1426
rect 13046 1392 13058 1426
rect 13058 1392 13080 1426
rect 13118 1392 13152 1426
rect 18994 2105 19100 2142
rect 18994 2071 19091 2105
rect 19091 2071 19100 2105
rect 18994 2034 19100 2071
rect 18994 2000 19091 2034
rect 19091 2000 19100 2034
rect 18994 1963 19100 2000
rect 18994 1929 19091 1963
rect 19091 1929 19100 1963
rect 18994 1892 19100 1929
rect 18994 1858 19091 1892
rect 19091 1858 19100 1892
rect 18994 1821 19100 1858
rect 18994 1787 19091 1821
rect 19091 1787 19100 1821
rect 18994 1750 19100 1787
rect 18994 1716 19091 1750
rect 19091 1716 19100 1750
rect 18994 1679 19100 1716
rect 18994 1645 19091 1679
rect 19091 1645 19100 1679
rect 18994 1608 19100 1645
rect 18994 1574 19091 1608
rect 19091 1574 19100 1608
rect 18994 1537 19100 1574
rect 18994 1503 19091 1537
rect 19091 1503 19100 1537
rect 18994 1466 19100 1503
rect 18994 1432 19091 1466
rect 19091 1432 19100 1466
rect 18994 1396 19100 1432
rect 10619 1282 10653 1316
rect 10619 1210 10653 1244
rect 10619 1138 10653 1172
rect 10619 1066 10653 1100
rect 10619 994 10653 1028
rect 10619 922 10653 956
rect 18994 1362 19091 1396
rect 19091 1362 19100 1396
rect 18994 1326 19100 1362
rect 18994 1301 19091 1326
rect 19091 1301 19100 1326
rect 18994 1228 19028 1262
rect 19066 1256 19100 1262
rect 19066 1228 19091 1256
rect 19091 1228 19100 1256
rect 18994 1155 19028 1189
rect 19066 1186 19100 1189
rect 19066 1155 19091 1186
rect 19091 1155 19100 1186
rect 18994 1082 19028 1116
rect 19066 1082 19091 1116
rect 19091 1082 19100 1116
rect 18994 1009 19028 1043
rect 19066 1012 19091 1043
rect 19091 1012 19100 1043
rect 19066 1009 19100 1012
rect 18994 936 19028 970
rect 19066 942 19091 970
rect 19091 942 19100 970
rect 19066 936 19100 942
rect 10619 850 10653 884
rect 10619 778 10653 812
rect 10619 706 10653 740
rect 10619 634 10653 668
rect 10619 562 10653 596
rect 10619 490 10653 524
rect 10619 428 10653 452
rect 19114 703 19148 737
rect 19114 622 19148 656
rect 19114 541 19148 575
rect 19114 460 19148 494
rect 10619 418 10653 428
rect 10619 346 10653 380
rect 19114 379 19148 413
rect 10619 304 10653 308
rect 10619 274 10653 304
rect 10619 214 10653 235
rect 10619 201 10653 214
rect 10619 158 10653 162
rect 10619 128 10653 158
rect 19114 298 19148 332
rect 19114 217 19148 251
rect 10729 90 10755 124
rect 10755 90 10763 124
rect 10801 90 10823 124
rect 10823 90 10835 124
rect 10873 90 10891 124
rect 10891 90 10907 124
rect 10945 90 10959 124
rect 10959 90 10979 124
rect 11017 90 11027 124
rect 11027 90 11051 124
rect 11089 90 11095 124
rect 11095 90 11123 124
rect 11161 90 11163 124
rect 11163 90 11195 124
rect 11233 90 11265 124
rect 11265 90 11267 124
rect 11305 90 11333 124
rect 11333 90 11339 124
rect 11377 90 11401 124
rect 11401 90 11411 124
rect 11449 90 11469 124
rect 11469 90 11483 124
rect 11521 90 11537 124
rect 11537 90 11555 124
rect 11593 90 11605 124
rect 11605 90 11627 124
rect 11665 90 11673 124
rect 11673 90 11699 124
rect 11737 90 11741 124
rect 11741 90 11771 124
rect 11809 90 11843 124
rect 11881 90 11911 124
rect 11911 90 11915 124
rect 11953 90 11979 124
rect 11979 90 11987 124
rect 12025 90 12047 124
rect 12047 90 12059 124
rect 12097 90 12115 124
rect 12115 90 12131 124
rect 12169 90 12183 124
rect 12183 90 12203 124
rect 12241 90 12251 124
rect 12251 90 12275 124
rect 12313 90 12319 124
rect 12319 90 12347 124
rect 12385 90 12387 124
rect 12387 90 12419 124
rect 12457 90 12489 124
rect 12489 90 12491 124
rect 12529 90 12557 124
rect 12557 90 12563 124
rect 12601 90 12625 124
rect 12625 90 12635 124
rect 12673 90 12693 124
rect 12693 90 12707 124
rect 12745 90 12761 124
rect 12761 90 12779 124
rect 12817 90 12829 124
rect 12829 90 12851 124
rect 12889 90 12897 124
rect 12897 90 12923 124
rect 12961 90 12965 124
rect 12965 90 12995 124
rect 13033 90 13067 124
rect 13105 90 13139 124
rect 13177 90 13211 124
rect 13249 90 13283 124
rect 13321 90 13355 124
rect 13393 90 13427 124
rect 13465 90 13499 124
rect 13537 90 13571 124
rect 13609 90 13643 124
rect 13681 90 13715 124
rect 13753 90 13787 124
rect 13825 90 13859 124
rect 13897 90 13931 124
rect 13969 90 14003 124
rect 14041 90 14075 124
rect 14113 90 14147 124
rect 14185 90 14219 124
rect 14258 90 14292 124
rect 14331 90 14365 124
rect 14404 90 14438 124
rect 14477 90 14511 124
rect 14550 90 14584 124
rect 14623 90 14657 124
rect 14696 90 14730 124
rect 14769 90 14803 124
rect 14842 90 14876 124
rect 14915 90 14949 124
rect 14988 90 15022 124
rect 15061 90 15095 124
rect 15134 90 15141 124
rect 15141 90 15168 124
rect 15207 90 15209 124
rect 15209 90 15241 124
rect 15280 90 15311 124
rect 15311 90 15314 124
rect 15353 90 15379 124
rect 15379 90 15387 124
rect 15426 90 15447 124
rect 15447 90 15460 124
rect 15499 90 15515 124
rect 15515 90 15533 124
rect 15572 90 15583 124
rect 15583 90 15606 124
rect 15645 90 15651 124
rect 15651 90 15679 124
rect 15718 90 15719 124
rect 15719 90 15752 124
rect 15791 90 15821 124
rect 15821 90 15825 124
rect 15864 90 15889 124
rect 15889 90 15898 124
rect 15937 90 15957 124
rect 15957 90 15971 124
rect 16010 90 16025 124
rect 16025 90 16044 124
rect 16083 90 16093 124
rect 16093 90 16117 124
rect 16156 90 16161 124
rect 16161 90 16190 124
rect 16229 90 16263 124
rect 16302 90 16331 124
rect 16331 90 16336 124
rect 16375 90 16399 124
rect 16399 90 16409 124
rect 16448 90 16467 124
rect 16467 90 16482 124
rect 16521 90 16535 124
rect 16535 90 16555 124
rect 16594 90 16603 124
rect 16603 90 16628 124
rect 16667 90 16671 124
rect 16671 90 16701 124
rect 16740 90 16773 124
rect 16773 90 16774 124
rect 16813 90 16841 124
rect 16841 90 16847 124
rect 16886 90 16909 124
rect 16909 90 16920 124
rect 16959 90 16977 124
rect 16977 90 16993 124
rect 17032 90 17045 124
rect 17045 90 17066 124
rect 17105 90 17113 124
rect 17113 90 17139 124
rect 17178 90 17181 124
rect 17181 90 17212 124
rect 17251 90 17283 124
rect 17283 90 17285 124
rect 17324 90 17351 124
rect 17351 90 17358 124
rect 17397 90 17419 124
rect 17419 90 17431 124
rect 17470 90 17487 124
rect 17487 90 17504 124
rect 17543 90 17555 124
rect 17555 90 17577 124
rect 17616 90 17623 124
rect 17623 90 17650 124
rect 17689 90 17691 124
rect 17691 90 17723 124
rect 17762 90 17793 124
rect 17793 90 17796 124
rect 17835 90 17861 124
rect 17861 90 17869 124
rect 17908 90 17929 124
rect 17929 90 17942 124
rect 17981 90 17997 124
rect 17997 90 18015 124
rect 18054 90 18065 124
rect 18065 90 18088 124
rect 18127 90 18133 124
rect 18133 90 18161 124
rect 18200 90 18201 124
rect 18201 90 18234 124
rect 18273 90 18303 124
rect 18303 90 18307 124
rect 18346 90 18371 124
rect 18371 90 18380 124
rect 18419 90 18439 124
rect 18439 90 18453 124
rect 18492 90 18507 124
rect 18507 90 18526 124
rect 18565 90 18575 124
rect 18575 90 18599 124
rect 18638 90 18643 124
rect 18643 90 18672 124
rect 18711 90 18745 124
rect 18784 90 18813 124
rect 18813 90 18818 124
rect 18857 90 18881 124
rect 18881 90 18891 124
rect 18930 90 18949 124
rect 18949 90 18964 124
rect 19003 90 19018 124
rect 19018 90 19037 124
rect 19076 90 19110 124
<< metal1 >>
rect 853 6908 13367 6914
rect 853 6874 865 6908
rect 899 6874 938 6908
rect 972 6874 1011 6908
rect 1045 6874 1084 6908
rect 1118 6874 1157 6908
rect 1191 6874 1230 6908
rect 1264 6874 1303 6908
rect 1337 6874 1376 6908
rect 1410 6874 1449 6908
rect 1483 6874 1522 6908
rect 1556 6874 1595 6908
rect 1629 6874 1668 6908
rect 1702 6874 1741 6908
rect 1775 6874 1814 6908
rect 1848 6874 1887 6908
rect 1921 6874 1960 6908
rect 1994 6874 2033 6908
rect 2067 6874 2106 6908
rect 2140 6874 2179 6908
rect 2213 6874 2252 6908
rect 853 6836 2252 6874
rect 853 6802 865 6836
rect 899 6802 938 6836
rect 972 6802 1011 6836
rect 1045 6802 1084 6836
rect 1118 6802 1157 6836
rect 1191 6802 1230 6836
rect 1264 6802 1303 6836
rect 1337 6802 1376 6836
rect 1410 6802 1449 6836
rect 1483 6802 1522 6836
rect 1556 6802 1595 6836
rect 1629 6802 1668 6836
rect 1702 6802 1741 6836
rect 1775 6802 1814 6836
rect 1848 6802 1887 6836
rect 1921 6802 1960 6836
rect 1994 6802 2033 6836
rect 2067 6802 2106 6836
rect 2140 6802 2179 6836
rect 2213 6802 2252 6836
rect 853 6796 13197 6802
tri 5716 6730 5782 6796 ne
rect 5782 6730 6515 6796
tri 6515 6730 6581 6796 nw
tri 13165 6771 13190 6796 ne
rect 13190 6730 13197 6796
rect 13302 6764 13367 6908
rect 13303 6730 13367 6764
tri 5782 6691 5821 6730 ne
rect 5821 6691 6476 6730
tri 6476 6691 6515 6730 nw
rect 13190 6691 13367 6730
tri 5821 6667 5845 6691 ne
rect 5845 6667 6442 6691
tri 5845 6654 5858 6667 ne
rect 5858 6633 5870 6667
rect 5904 6633 5945 6667
rect 5979 6633 6020 6667
rect 6054 6633 6095 6667
rect 6129 6633 6170 6667
rect 6204 6633 6245 6667
rect 6279 6633 6319 6667
rect 6353 6633 6393 6667
rect 6427 6657 6442 6667
tri 6442 6657 6476 6691 nw
rect 13190 6657 13197 6691
rect 13231 6657 13269 6691
rect 13303 6657 13367 6691
rect 6427 6633 6439 6657
tri 6439 6654 6442 6657 nw
rect 5858 6627 6439 6633
rect 13190 6618 13367 6657
rect 13190 6584 13197 6618
rect 13231 6584 13269 6618
rect 13303 6584 13367 6618
rect 5786 6563 6452 6575
rect 5786 6529 5792 6563
rect 5826 6529 6452 6563
rect 5786 6523 6452 6529
rect 6504 6523 6516 6575
rect 6568 6523 6574 6575
rect 5786 6491 5832 6523
tri 5832 6498 5857 6523 nw
tri 6491 6498 6516 6523 ne
rect 5786 6457 5792 6491
rect 5826 6457 5832 6491
rect 5786 6445 5832 6457
rect 6516 6491 6562 6523
tri 6562 6511 6574 6523 nw
rect 13190 6545 13367 6584
rect 6516 6457 6522 6491
rect 6556 6457 6562 6491
rect 6516 6445 6562 6457
rect 5858 6411 6560 6417
rect 5858 6377 5870 6411
rect 5904 6377 5945 6411
rect 5979 6377 6020 6411
rect 6054 6377 6095 6411
rect 6129 6377 6170 6411
rect 6204 6377 6245 6411
rect 6279 6377 6319 6411
rect 6353 6377 6393 6411
rect 6427 6377 6560 6411
rect 5858 6301 6560 6377
rect 6561 6302 6562 6416
rect 6598 6302 6599 6416
rect 6600 6301 6625 6417
rect 6805 6301 6811 6417
tri 6846 6378 6880 6412 se
rect 6880 6378 13111 6412
rect 6846 6366 13111 6378
rect 6846 6338 6892 6366
tri 6892 6341 6917 6366 nw
tri 13091 6346 13111 6366 ne
tri 13111 6361 13162 6412 sw
rect 13111 6346 13162 6361
tri 13111 6341 13116 6346 ne
rect 6847 6336 6891 6337
rect 6846 6300 6892 6336
rect 6847 6299 6891 6300
rect 6846 6281 6892 6298
rect 6846 6247 6852 6281
rect 6886 6247 6892 6281
rect 6846 6209 6892 6247
rect 6846 6175 6852 6209
rect 6886 6175 6892 6209
rect 6846 6081 6892 6175
rect 6847 6079 6891 6080
rect 6846 6043 6892 6079
rect 6847 6042 6891 6043
rect 6846 5931 6892 6041
rect 6846 5897 6852 5931
rect 6886 5897 6892 5931
rect 6846 5859 6892 5897
rect 6846 5825 6852 5859
rect 6886 5825 6892 5859
rect 6846 5645 6892 5825
rect 6847 5643 6891 5644
rect 6846 5613 6892 5643
rect 6847 5612 6891 5613
rect 6846 5584 6892 5611
rect 6846 5550 6852 5584
rect 6886 5550 6892 5584
rect 6846 5512 6892 5550
rect 6846 5478 6852 5512
rect 6886 5478 6892 5512
rect 6846 5309 6892 5478
rect 6847 5307 6891 5308
rect 6846 5277 6892 5307
rect 6847 5276 6891 5277
rect 6846 5244 6892 5275
rect 6846 5210 6852 5244
rect 6886 5210 6892 5244
rect 6920 6323 9892 6329
rect 6920 6289 6932 6323
rect 6966 6289 7005 6323
rect 7039 6289 7078 6323
rect 7112 6289 7151 6323
rect 7185 6289 7224 6323
rect 7258 6289 7297 6323
rect 7331 6289 7370 6323
rect 7404 6289 7443 6323
rect 7477 6289 7516 6323
rect 7550 6289 7589 6323
rect 7623 6289 7662 6323
rect 7696 6289 7735 6323
rect 7769 6289 7808 6323
rect 7842 6289 7881 6323
rect 7915 6289 7954 6323
rect 7988 6289 8027 6323
rect 8061 6289 8100 6323
rect 8134 6289 8173 6323
rect 8207 6289 8246 6323
rect 8280 6289 8319 6323
rect 8353 6289 8392 6323
rect 8426 6289 8465 6323
rect 8499 6289 8538 6323
rect 8572 6289 8611 6323
rect 8645 6289 8684 6323
rect 8718 6289 8757 6323
rect 8791 6289 8830 6323
rect 8864 6289 8903 6323
rect 8937 6289 8976 6323
rect 9010 6289 9049 6323
rect 9083 6289 9122 6323
rect 9156 6289 9195 6323
rect 9229 6289 9268 6323
rect 9302 6289 9341 6323
rect 9375 6289 9414 6323
rect 9448 6289 9486 6323
rect 9520 6289 9558 6323
rect 9592 6289 9630 6323
rect 9664 6289 9702 6323
rect 9736 6289 9774 6323
rect 9808 6289 9846 6323
rect 9880 6289 9892 6323
rect 6920 6283 9892 6289
rect 10119 6323 13088 6329
rect 10119 6289 10131 6323
rect 10165 6289 10203 6323
rect 10237 6289 10275 6323
rect 10309 6289 10347 6323
rect 10381 6289 10419 6323
rect 10453 6289 10491 6323
rect 10525 6289 10563 6323
rect 10597 6289 10635 6323
rect 10669 6289 10707 6323
rect 10741 6289 10779 6323
rect 10813 6289 10852 6323
rect 10886 6289 10925 6323
rect 10959 6289 10998 6323
rect 11032 6289 11071 6323
rect 11105 6289 11144 6323
rect 11178 6289 11217 6323
rect 11251 6289 11290 6323
rect 11324 6289 11363 6323
rect 11397 6289 11436 6323
rect 11470 6289 11509 6323
rect 11543 6289 11582 6323
rect 11616 6289 11655 6323
rect 11689 6289 11728 6323
rect 11762 6289 11801 6323
rect 11835 6289 11874 6323
rect 11908 6289 11947 6323
rect 11981 6289 12020 6323
rect 12054 6289 12093 6323
rect 12127 6289 12166 6323
rect 12200 6289 12239 6323
rect 12273 6289 12312 6323
rect 12346 6289 12385 6323
rect 12419 6289 12458 6323
rect 12492 6289 12531 6323
rect 12565 6289 12604 6323
rect 12638 6289 12677 6323
rect 12711 6289 12750 6323
rect 12784 6289 12823 6323
rect 12857 6289 12896 6323
rect 12930 6289 12969 6323
rect 13003 6289 13042 6323
rect 13076 6289 13088 6323
rect 10119 6283 13088 6289
rect 6920 6281 7155 6283
tri 7155 6281 7157 6283 nw
tri 12851 6281 12853 6283 ne
rect 12853 6281 13088 6283
rect 6920 5981 7132 6281
tri 7132 6258 7155 6281 nw
tri 12853 6258 12876 6281 ne
rect 7160 6167 9856 6173
rect 9858 6172 9894 6173
rect 7160 6133 7172 6167
rect 7206 6133 7246 6167
rect 7280 6133 7320 6167
rect 7354 6133 7394 6167
rect 7428 6133 7468 6167
rect 7502 6133 7542 6167
rect 7576 6133 7616 6167
rect 7650 6133 7690 6167
rect 7724 6133 7764 6167
rect 7798 6133 7837 6167
rect 7871 6133 7910 6167
rect 7944 6133 7983 6167
rect 8017 6133 8056 6167
rect 8090 6133 8129 6167
rect 8163 6133 8202 6167
rect 8236 6133 8275 6167
rect 8309 6133 8348 6167
rect 8382 6133 8421 6167
rect 8455 6133 8494 6167
rect 8528 6133 8567 6167
rect 8601 6133 8640 6167
rect 8674 6133 8713 6167
rect 8747 6133 8786 6167
rect 8820 6133 8859 6167
rect 8893 6133 8932 6167
rect 8966 6133 9005 6167
rect 9039 6133 9078 6167
rect 9112 6133 9151 6167
rect 9185 6133 9224 6167
rect 9258 6133 9297 6167
rect 9331 6133 9370 6167
rect 9404 6133 9443 6167
rect 9477 6133 9516 6167
rect 9550 6133 9589 6167
rect 9623 6133 9662 6167
rect 9696 6133 9735 6167
rect 9769 6133 9808 6167
rect 9842 6133 9856 6167
rect 7160 6127 9856 6133
rect 9857 6128 9895 6172
rect 9858 6127 9894 6128
rect 9896 6127 9989 6173
tri 9895 6102 9920 6127 ne
tri 7132 5981 7157 6006 sw
rect 6920 5975 9892 5981
rect 6920 5941 6932 5975
rect 6966 5941 7005 5975
rect 7039 5941 7078 5975
rect 7112 5941 7151 5975
rect 7185 5941 7224 5975
rect 7258 5941 7297 5975
rect 7331 5941 7370 5975
rect 7404 5941 7443 5975
rect 7477 5941 7516 5975
rect 7550 5941 7589 5975
rect 7623 5941 7662 5975
rect 7696 5941 7735 5975
rect 7769 5941 7808 5975
rect 7842 5941 7881 5975
rect 7915 5941 7954 5975
rect 7988 5941 8027 5975
rect 8061 5941 8100 5975
rect 8134 5941 8173 5975
rect 8207 5941 8246 5975
rect 8280 5941 8319 5975
rect 8353 5941 8392 5975
rect 8426 5941 8465 5975
rect 8499 5941 8538 5975
rect 8572 5941 8611 5975
rect 8645 5941 8684 5975
rect 8718 5941 8757 5975
rect 8791 5941 8830 5975
rect 8864 5941 8903 5975
rect 8937 5941 8976 5975
rect 9010 5941 9049 5975
rect 9083 5941 9122 5975
rect 9156 5941 9195 5975
rect 9229 5941 9268 5975
rect 9302 5941 9341 5975
rect 9375 5941 9414 5975
rect 9448 5941 9486 5975
rect 9520 5941 9558 5975
rect 9592 5941 9630 5975
rect 9664 5941 9702 5975
rect 9736 5941 9774 5975
rect 9808 5941 9846 5975
rect 9880 5941 9892 5975
rect 6920 5935 9892 5941
rect 6920 5933 7155 5935
tri 7155 5933 7157 5935 nw
rect 6920 5633 7132 5933
tri 7132 5910 7155 5933 nw
tri 9897 5827 9920 5850 se
rect 9920 5827 9989 6127
tri 9895 5825 9897 5827 se
rect 9897 5825 9989 5827
rect 7169 5819 9856 5825
rect 9858 5824 9894 5825
rect 7169 5785 7181 5819
rect 7215 5785 7254 5819
rect 7288 5785 7327 5819
rect 7361 5785 7400 5819
rect 7434 5785 7473 5819
rect 7507 5785 7546 5819
rect 7580 5785 7619 5819
rect 7653 5785 7692 5819
rect 7726 5785 7765 5819
rect 7799 5785 7838 5819
rect 7872 5785 7911 5819
rect 7945 5785 7984 5819
rect 8018 5785 8057 5819
rect 8091 5785 8130 5819
rect 8164 5785 8203 5819
rect 8237 5785 8276 5819
rect 8310 5785 8349 5819
rect 8383 5785 8422 5819
rect 8456 5785 8494 5819
rect 8528 5785 8566 5819
rect 8600 5785 8638 5819
rect 8672 5785 8710 5819
rect 8744 5785 8782 5819
rect 8816 5785 8854 5819
rect 8888 5785 8926 5819
rect 8960 5785 8998 5819
rect 9032 5785 9070 5819
rect 9104 5785 9142 5819
rect 9176 5785 9214 5819
rect 9248 5785 9286 5819
rect 9320 5785 9358 5819
rect 9392 5785 9430 5819
rect 9464 5785 9502 5819
rect 9536 5785 9574 5819
rect 9608 5785 9856 5819
rect 7169 5779 9856 5785
rect 9857 5780 9895 5824
rect 9858 5779 9894 5780
rect 9896 5779 9989 5825
tri 9895 5754 9920 5779 ne
tri 7132 5633 7157 5658 sw
rect 6920 5627 9892 5633
rect 6920 5593 6932 5627
rect 6966 5593 7005 5627
rect 7039 5593 7078 5627
rect 7112 5593 7151 5627
rect 7185 5593 7224 5627
rect 7258 5593 7297 5627
rect 7331 5593 7370 5627
rect 7404 5593 7443 5627
rect 7477 5593 7516 5627
rect 7550 5593 7589 5627
rect 7623 5593 7662 5627
rect 7696 5593 7735 5627
rect 7769 5593 7808 5627
rect 7842 5593 7881 5627
rect 7915 5593 7954 5627
rect 7988 5593 8027 5627
rect 8061 5593 8100 5627
rect 8134 5593 8173 5627
rect 8207 5593 8246 5627
rect 8280 5593 8319 5627
rect 8353 5593 8392 5627
rect 8426 5593 8465 5627
rect 8499 5593 8538 5627
rect 8572 5593 8611 5627
rect 8645 5593 8684 5627
rect 8718 5593 8757 5627
rect 8791 5593 8830 5627
rect 8864 5593 8903 5627
rect 8937 5593 8976 5627
rect 9010 5593 9049 5627
rect 9083 5593 9122 5627
rect 9156 5593 9195 5627
rect 9229 5593 9268 5627
rect 9302 5593 9341 5627
rect 9375 5593 9414 5627
rect 9448 5593 9486 5627
rect 9520 5593 9558 5627
rect 9592 5593 9630 5627
rect 9664 5593 9702 5627
rect 9736 5593 9774 5627
rect 9808 5593 9846 5627
rect 9880 5593 9892 5627
rect 6920 5587 9892 5593
rect 6920 5585 7155 5587
tri 7155 5585 7157 5587 nw
rect 6920 5285 7132 5585
tri 7132 5562 7155 5585 nw
tri 9897 5479 9920 5502 se
rect 9920 5479 9989 5779
tri 9895 5477 9897 5479 se
rect 9897 5477 9989 5479
rect 7160 5471 9856 5477
rect 9858 5476 9894 5477
rect 7160 5437 7172 5471
rect 7206 5437 7246 5471
rect 7280 5437 7320 5471
rect 7354 5437 7394 5471
rect 7428 5437 7468 5471
rect 7502 5437 7542 5471
rect 7576 5437 7616 5471
rect 7650 5437 7690 5471
rect 7724 5437 7764 5471
rect 7798 5437 7838 5471
rect 7872 5437 7912 5471
rect 7946 5437 7985 5471
rect 8019 5437 8058 5471
rect 8092 5437 8131 5471
rect 8165 5437 8204 5471
rect 8238 5437 8277 5471
rect 8311 5437 8350 5471
rect 8384 5437 8423 5471
rect 8457 5437 8496 5471
rect 8530 5437 8569 5471
rect 8603 5437 8642 5471
rect 8676 5437 8715 5471
rect 8749 5437 8788 5471
rect 8822 5437 8861 5471
rect 8895 5437 8934 5471
rect 8968 5437 9007 5471
rect 9041 5437 9080 5471
rect 9114 5437 9153 5471
rect 9187 5437 9226 5471
rect 9260 5437 9299 5471
rect 9333 5437 9372 5471
rect 9406 5437 9445 5471
rect 9479 5437 9518 5471
rect 9552 5437 9591 5471
rect 9625 5437 9664 5471
rect 9698 5437 9737 5471
rect 9771 5437 9810 5471
rect 9844 5437 9856 5471
rect 7160 5431 9856 5437
rect 9857 5432 9895 5476
rect 9858 5431 9894 5432
rect 9896 5431 9989 5477
tri 9895 5406 9920 5431 ne
tri 7132 5285 7157 5310 sw
rect 6920 5279 9892 5285
rect 6920 5245 6932 5279
rect 6966 5245 7005 5279
rect 7039 5245 7078 5279
rect 7112 5245 7151 5279
rect 7185 5245 7224 5279
rect 7258 5245 7297 5279
rect 7331 5245 7370 5279
rect 7404 5245 7443 5279
rect 7477 5245 7516 5279
rect 7550 5245 7589 5279
rect 7623 5245 7662 5279
rect 7696 5245 7735 5279
rect 7769 5245 7808 5279
rect 7842 5245 7881 5279
rect 7915 5245 7954 5279
rect 7988 5245 8027 5279
rect 8061 5245 8100 5279
rect 8134 5245 8173 5279
rect 8207 5245 8246 5279
rect 8280 5245 8319 5279
rect 8353 5245 8392 5279
rect 8426 5245 8465 5279
rect 8499 5245 8538 5279
rect 8572 5245 8611 5279
rect 8645 5245 8684 5279
rect 8718 5245 8757 5279
rect 8791 5245 8830 5279
rect 8864 5245 8903 5279
rect 8937 5245 8976 5279
rect 9010 5245 9049 5279
rect 9083 5245 9122 5279
rect 9156 5245 9195 5279
rect 9229 5245 9268 5279
rect 9302 5245 9341 5279
rect 9375 5245 9414 5279
rect 9448 5245 9486 5279
rect 9520 5245 9558 5279
rect 9592 5245 9630 5279
rect 9664 5245 9702 5279
rect 9736 5245 9774 5279
rect 9808 5245 9846 5279
rect 9880 5245 9892 5279
rect 6920 5239 9892 5245
tri 6829 5180 6846 5197 se
rect 6846 5180 6892 5210
tri 6821 5172 6829 5180 se
rect 6829 5172 6892 5180
rect 6696 5126 6780 5172
rect 6781 5127 6782 5171
rect 6812 5127 6813 5171
rect 6814 5138 6852 5172
rect 6886 5138 6892 5172
rect 6814 5126 6892 5138
rect 6920 5123 9833 5129
rect 6920 5089 6932 5123
rect 6966 5089 7006 5123
rect 7040 5089 7080 5123
rect 7114 5089 7154 5123
rect 7188 5089 7228 5123
rect 7262 5089 7302 5123
rect 7336 5089 7376 5123
rect 7410 5089 7450 5123
rect 7484 5089 7524 5123
rect 7558 5089 7597 5123
rect 7631 5089 7670 5123
rect 7704 5089 7743 5123
rect 7777 5089 7816 5123
rect 7850 5089 7889 5123
rect 7923 5089 7962 5123
rect 7996 5089 8035 5123
rect 8069 5089 8108 5123
rect 8142 5089 8181 5123
rect 8215 5089 8254 5123
rect 8288 5089 8327 5123
rect 8361 5089 8400 5123
rect 8434 5089 8473 5123
rect 8507 5089 8546 5123
rect 8580 5089 8619 5123
rect 8653 5089 8692 5123
rect 8726 5089 8765 5123
rect 8799 5089 8838 5123
rect 8872 5089 8911 5123
rect 8945 5089 8984 5123
rect 9018 5089 9057 5123
rect 9091 5089 9130 5123
rect 9164 5089 9203 5123
rect 9237 5089 9276 5123
rect 9310 5089 9349 5123
rect 9383 5089 9422 5123
rect 9456 5089 9495 5123
rect 9529 5089 9568 5123
rect 9602 5089 9641 5123
rect 9675 5089 9714 5123
rect 9748 5089 9787 5123
rect 9821 5089 9833 5123
rect 6920 5085 9833 5089
rect 6921 5083 9832 5084
rect 6920 5055 9833 5083
rect 6921 5054 9832 5055
tri 6905 5039 6920 5054 se
tri 9833 5053 9834 5054 sw
tri 9919 5053 9920 5054 se
rect 9920 5053 9989 5431
rect 6920 5039 9834 5053
tri 6811 5029 6821 5039 sw
tri 6895 5029 6905 5039 se
rect 6905 5029 9834 5039
tri 9834 5029 9858 5053 sw
tri 9895 5029 9919 5053 se
rect 9919 5029 9989 5053
rect 6811 4859 9989 5029
rect 10021 6127 10115 6173
rect 10117 6172 10153 6173
rect 10116 6128 10154 6172
rect 10155 6167 12848 6173
rect 10155 6133 10169 6167
rect 10203 6133 10242 6167
rect 10276 6133 10315 6167
rect 10349 6133 10388 6167
rect 10422 6133 10461 6167
rect 10495 6133 10534 6167
rect 10568 6133 10607 6167
rect 10641 6133 10680 6167
rect 10714 6133 10753 6167
rect 10787 6133 10826 6167
rect 10860 6133 10899 6167
rect 10933 6133 10972 6167
rect 11006 6133 11045 6167
rect 11079 6133 11118 6167
rect 11152 6133 11191 6167
rect 11225 6133 11264 6167
rect 11298 6133 11337 6167
rect 11371 6133 11410 6167
rect 11444 6133 11483 6167
rect 11517 6133 11556 6167
rect 11590 6133 11629 6167
rect 11663 6133 11702 6167
rect 11736 6133 11775 6167
rect 11809 6133 11848 6167
rect 11882 6133 11921 6167
rect 11955 6133 11994 6167
rect 12028 6133 12067 6167
rect 12101 6133 12140 6167
rect 12174 6133 12213 6167
rect 12247 6133 12286 6167
rect 12320 6133 12359 6167
rect 12393 6133 12432 6167
rect 12466 6133 12506 6167
rect 12540 6133 12580 6167
rect 12614 6133 12654 6167
rect 12688 6133 12728 6167
rect 12762 6133 12802 6167
rect 12836 6133 12848 6167
rect 10117 6127 10153 6128
rect 10155 6127 12848 6133
rect 10021 5827 10091 6127
tri 10091 6102 10116 6127 nw
tri 12851 5981 12876 6006 se
rect 12876 5981 13088 6281
rect 10119 5975 13088 5981
rect 10119 5941 10131 5975
rect 10165 5941 10203 5975
rect 10237 5941 10275 5975
rect 10309 5941 10347 5975
rect 10381 5941 10419 5975
rect 10453 5941 10491 5975
rect 10525 5941 10563 5975
rect 10597 5941 10635 5975
rect 10669 5941 10707 5975
rect 10741 5941 10779 5975
rect 10813 5941 10852 5975
rect 10886 5941 10925 5975
rect 10959 5941 10998 5975
rect 11032 5941 11071 5975
rect 11105 5941 11144 5975
rect 11178 5941 11217 5975
rect 11251 5941 11290 5975
rect 11324 5941 11363 5975
rect 11397 5941 11436 5975
rect 11470 5941 11509 5975
rect 11543 5941 11582 5975
rect 11616 5941 11655 5975
rect 11689 5941 11728 5975
rect 11762 5941 11801 5975
rect 11835 5941 11874 5975
rect 11908 5941 11947 5975
rect 11981 5941 12020 5975
rect 12054 5941 12093 5975
rect 12127 5941 12166 5975
rect 12200 5941 12239 5975
rect 12273 5941 12312 5975
rect 12346 5941 12385 5975
rect 12419 5941 12458 5975
rect 12492 5941 12531 5975
rect 12565 5941 12604 5975
rect 12638 5941 12677 5975
rect 12711 5941 12750 5975
rect 12784 5941 12823 5975
rect 12857 5941 12896 5975
rect 12930 5941 12969 5975
rect 13003 5941 13042 5975
rect 13076 5941 13088 5975
rect 10119 5935 13088 5941
tri 12851 5933 12853 5935 ne
rect 12853 5933 13088 5935
tri 12853 5910 12876 5933 ne
tri 10091 5827 10114 5850 sw
rect 10021 5825 10114 5827
tri 10114 5825 10116 5827 sw
rect 10021 5779 10115 5825
rect 10117 5824 10153 5825
rect 10116 5780 10154 5824
rect 10155 5819 12848 5825
rect 10155 5785 10169 5819
rect 10203 5785 10242 5819
rect 10276 5785 10315 5819
rect 10349 5785 10388 5819
rect 10422 5785 10461 5819
rect 10495 5785 10534 5819
rect 10568 5785 10607 5819
rect 10641 5785 10680 5819
rect 10714 5785 10753 5819
rect 10787 5785 10826 5819
rect 10860 5785 10899 5819
rect 10933 5785 10972 5819
rect 11006 5785 11045 5819
rect 11079 5785 11118 5819
rect 11152 5785 11191 5819
rect 11225 5785 11264 5819
rect 11298 5785 11337 5819
rect 11371 5785 11410 5819
rect 11444 5785 11483 5819
rect 11517 5785 11556 5819
rect 11590 5785 11629 5819
rect 11663 5785 11702 5819
rect 11736 5785 11775 5819
rect 11809 5785 11848 5819
rect 11882 5785 11921 5819
rect 11955 5785 11994 5819
rect 12028 5785 12067 5819
rect 12101 5785 12140 5819
rect 12174 5785 12213 5819
rect 12247 5785 12286 5819
rect 12320 5785 12359 5819
rect 12393 5785 12432 5819
rect 12466 5785 12506 5819
rect 12540 5785 12580 5819
rect 12614 5785 12654 5819
rect 12688 5785 12728 5819
rect 12762 5785 12802 5819
rect 12836 5785 12848 5819
rect 10117 5779 10153 5780
rect 10155 5779 12848 5785
rect 10021 5479 10091 5779
tri 10091 5754 10116 5779 nw
tri 12851 5633 12876 5658 se
rect 12876 5633 13088 5933
rect 10119 5627 13088 5633
rect 10119 5593 10131 5627
rect 10165 5593 10203 5627
rect 10237 5593 10275 5627
rect 10309 5593 10347 5627
rect 10381 5593 10419 5627
rect 10453 5593 10491 5627
rect 10525 5593 10563 5627
rect 10597 5593 10635 5627
rect 10669 5593 10707 5627
rect 10741 5593 10779 5627
rect 10813 5593 10852 5627
rect 10886 5593 10925 5627
rect 10959 5593 10998 5627
rect 11032 5593 11071 5627
rect 11105 5593 11144 5627
rect 11178 5593 11217 5627
rect 11251 5593 11290 5627
rect 11324 5593 11363 5627
rect 11397 5593 11436 5627
rect 11470 5593 11509 5627
rect 11543 5593 11582 5627
rect 11616 5593 11655 5627
rect 11689 5593 11728 5627
rect 11762 5593 11801 5627
rect 11835 5593 11874 5627
rect 11908 5593 11947 5627
rect 11981 5593 12020 5627
rect 12054 5593 12093 5627
rect 12127 5593 12166 5627
rect 12200 5593 12239 5627
rect 12273 5593 12312 5627
rect 12346 5593 12385 5627
rect 12419 5593 12458 5627
rect 12492 5593 12531 5627
rect 12565 5593 12604 5627
rect 12638 5593 12677 5627
rect 12711 5593 12750 5627
rect 12784 5593 12823 5627
rect 12857 5593 12896 5627
rect 12930 5593 12969 5627
rect 13003 5593 13042 5627
rect 13076 5593 13088 5627
rect 10119 5587 13088 5593
tri 12851 5585 12853 5587 ne
rect 12853 5585 13088 5587
tri 12853 5562 12876 5585 ne
tri 10091 5479 10114 5502 sw
rect 10021 5477 10114 5479
tri 10114 5477 10116 5479 sw
rect 10021 5431 10115 5477
rect 10117 5476 10153 5477
rect 10116 5432 10154 5476
rect 10155 5471 12848 5477
rect 10155 5437 10169 5471
rect 10203 5437 10242 5471
rect 10276 5437 10315 5471
rect 10349 5437 10388 5471
rect 10422 5437 10461 5471
rect 10495 5437 10534 5471
rect 10568 5437 10607 5471
rect 10641 5437 10680 5471
rect 10714 5437 10753 5471
rect 10787 5437 10826 5471
rect 10860 5437 10899 5471
rect 10933 5437 10972 5471
rect 11006 5437 11045 5471
rect 11079 5437 11118 5471
rect 11152 5437 11191 5471
rect 11225 5437 11264 5471
rect 11298 5437 11337 5471
rect 11371 5437 11410 5471
rect 11444 5437 11483 5471
rect 11517 5437 11556 5471
rect 11590 5437 11629 5471
rect 11663 5437 11702 5471
rect 11736 5437 11775 5471
rect 11809 5437 11848 5471
rect 11882 5437 11921 5471
rect 11955 5437 11994 5471
rect 12028 5437 12067 5471
rect 12101 5437 12140 5471
rect 12174 5437 12213 5471
rect 12247 5437 12286 5471
rect 12320 5437 12359 5471
rect 12393 5437 12432 5471
rect 12466 5437 12506 5471
rect 12540 5437 12580 5471
rect 12614 5437 12654 5471
rect 12688 5437 12728 5471
rect 12762 5437 12802 5471
rect 12836 5437 12848 5471
rect 10117 5431 10153 5432
rect 10155 5431 12848 5437
rect 10021 5029 10091 5431
tri 10091 5406 10116 5431 nw
tri 12851 5285 12876 5310 se
rect 12876 5285 13088 5585
rect 10119 5279 13088 5285
rect 10119 5245 10131 5279
rect 10165 5245 10203 5279
rect 10237 5245 10275 5279
rect 10309 5245 10347 5279
rect 10381 5245 10419 5279
rect 10453 5245 10491 5279
rect 10525 5245 10563 5279
rect 10597 5245 10635 5279
rect 10669 5245 10707 5279
rect 10741 5245 10779 5279
rect 10813 5245 10852 5279
rect 10886 5245 10925 5279
rect 10959 5245 10998 5279
rect 11032 5245 11071 5279
rect 11105 5245 11144 5279
rect 11178 5245 11217 5279
rect 11251 5245 11290 5279
rect 11324 5245 11363 5279
rect 11397 5245 11436 5279
rect 11470 5245 11509 5279
rect 11543 5245 11582 5279
rect 11616 5245 11655 5279
rect 11689 5245 11728 5279
rect 11762 5245 11801 5279
rect 11835 5245 11874 5279
rect 11908 5245 11947 5279
rect 11981 5245 12020 5279
rect 12054 5245 12093 5279
rect 12127 5245 12166 5279
rect 12200 5245 12239 5279
rect 12273 5245 12312 5279
rect 12346 5245 12385 5279
rect 12419 5245 12458 5279
rect 12492 5245 12531 5279
rect 12565 5245 12604 5279
rect 12638 5245 12677 5279
rect 12711 5245 12750 5279
rect 12784 5245 12823 5279
rect 12857 5245 12896 5279
rect 12930 5245 12969 5279
rect 13003 5245 13042 5279
rect 13076 5245 13088 5279
rect 10119 5239 13088 5245
rect 13116 6281 13162 6346
rect 13116 6247 13122 6281
rect 13156 6247 13162 6281
rect 13116 6209 13162 6247
rect 13116 6175 13122 6209
rect 13156 6175 13162 6209
rect 13116 6153 13162 6175
rect 13117 6151 13161 6152
rect 13116 6115 13162 6151
rect 13117 6114 13161 6115
rect 13116 5933 13162 6113
rect 13116 5899 13122 5933
rect 13156 5899 13162 5933
rect 13116 5861 13162 5899
rect 13116 5827 13122 5861
rect 13156 5827 13162 5861
rect 13116 5805 13162 5827
rect 13117 5803 13161 5804
rect 13116 5767 13162 5803
rect 13117 5766 13161 5767
rect 13116 5585 13162 5765
rect 13116 5551 13122 5585
rect 13156 5551 13162 5585
rect 13116 5513 13162 5551
rect 13116 5479 13122 5513
rect 13156 5479 13162 5513
rect 13116 5409 13162 5479
rect 13117 5407 13161 5408
rect 13116 5371 13162 5407
rect 13117 5370 13161 5371
rect 13116 5252 13162 5369
rect 13116 5218 13122 5252
rect 13156 5218 13162 5252
rect 13116 5180 13162 5218
rect 13116 5146 13122 5180
rect 13156 5146 13162 5180
rect 13116 5134 13162 5146
rect 13117 5132 13161 5133
rect 10184 5123 13088 5129
rect 10184 5089 10196 5123
rect 10230 5089 10268 5123
rect 10302 5089 10341 5123
rect 10375 5089 10414 5123
rect 10448 5089 10487 5123
rect 10521 5089 10560 5123
rect 10594 5089 10633 5123
rect 10667 5089 10706 5123
rect 10740 5089 10779 5123
rect 10813 5089 10852 5123
rect 10886 5089 10925 5123
rect 10959 5089 10998 5123
rect 11032 5089 11071 5123
rect 11105 5089 11144 5123
rect 11178 5089 11217 5123
rect 11251 5089 11290 5123
rect 11324 5089 11363 5123
rect 11397 5089 11436 5123
rect 11470 5089 11509 5123
rect 11543 5089 11582 5123
rect 11616 5089 11655 5123
rect 11689 5089 11728 5123
rect 11762 5089 11801 5123
rect 11835 5089 11874 5123
rect 11908 5089 11947 5123
rect 11981 5089 12020 5123
rect 12054 5089 12093 5123
rect 12127 5089 12166 5123
rect 12200 5089 12239 5123
rect 12273 5089 12312 5123
rect 12346 5089 12385 5123
rect 12419 5089 12458 5123
rect 12492 5089 12531 5123
rect 12565 5089 12604 5123
rect 12638 5089 12677 5123
rect 12711 5089 12750 5123
rect 12784 5089 12823 5123
rect 12857 5089 12896 5123
rect 12930 5089 12969 5123
rect 13003 5089 13042 5123
rect 13076 5089 13088 5123
rect 10184 5085 13088 5089
rect 10185 5083 13087 5084
rect 10184 5055 13088 5083
rect 13116 5096 13162 5132
rect 13190 5143 13197 6545
rect 13303 5143 13367 6545
rect 13190 5102 13367 5143
tri 13311 5096 13317 5102 ne
rect 13317 5096 13367 5102
rect 13117 5095 13161 5096
tri 13317 5095 13318 5096 ne
rect 13318 5095 13367 5096
tri 13318 5094 13319 5095 ne
rect 13319 5094 13367 5095
rect 13116 5081 13162 5094
tri 13319 5086 13327 5094 ne
rect 13327 5086 13367 5094
tri 13162 5081 13167 5086 sw
tri 13327 5081 13332 5086 ne
rect 13332 5081 13367 5086
rect 13116 5066 13167 5081
tri 13116 5055 13127 5066 ne
rect 13127 5061 13167 5066
tri 13167 5061 13187 5081 sw
tri 13332 5077 13336 5081 ne
rect 13127 5055 13267 5061
rect 10185 5054 13087 5055
tri 13127 5054 13128 5055 ne
rect 13128 5054 13267 5055
tri 10091 5029 10116 5054 sw
tri 10159 5029 10184 5054 se
tri 13088 5053 13089 5054 sw
tri 13128 5053 13129 5054 ne
rect 13129 5053 13267 5054
rect 10184 5029 13089 5053
rect 10021 5026 13089 5029
tri 13089 5026 13116 5053 sw
tri 13129 5026 13156 5053 ne
rect 13156 5026 13267 5053
rect 10021 5015 13116 5026
tri 13116 5015 13127 5026 sw
tri 13156 5015 13167 5026 ne
rect 13167 5020 13267 5026
tri 13267 5020 13308 5061 sw
rect 13167 5015 13308 5020
rect 10021 4975 13127 5015
tri 13127 4975 13167 5015 sw
tri 13240 4987 13268 5015 ne
rect 10021 4859 13118 4975
rect 13234 4859 13240 4975
tri 13243 4822 13268 4847 se
rect 13268 4822 13308 5015
rect 6770 4821 13308 4822
rect 6770 4817 13252 4821
rect 6770 4765 6776 4817
rect 6828 4765 6840 4817
rect 6892 4765 13252 4817
tri 13252 4765 13308 4821 nw
tri 13311 4737 13336 4762 se
rect 13336 4737 13367 5081
rect 3366 4731 13367 4737
rect 3366 4697 3410 4731
rect 3444 4697 3483 4731
rect 3517 4697 3556 4731
rect 3590 4697 3629 4731
rect 3663 4697 3702 4731
rect 3736 4697 3775 4731
rect 3809 4697 3848 4731
rect 3882 4697 3921 4731
rect 3955 4697 3994 4731
rect 4028 4697 4067 4731
rect 4101 4697 4140 4731
rect 4174 4697 4213 4731
rect 4247 4697 4286 4731
rect 4320 4697 4359 4731
rect 4393 4697 4432 4731
rect 4466 4697 4505 4731
rect 4539 4697 4578 4731
rect 4612 4697 4651 4731
rect 4685 4697 4724 4731
rect 4758 4697 4797 4731
rect 4831 4697 4870 4731
rect 4904 4697 4943 4731
rect 4977 4697 5016 4731
rect 5050 4697 5089 4731
rect 5123 4697 5162 4731
rect 5196 4697 5235 4731
rect 5269 4697 5307 4731
rect 5341 4697 5379 4731
rect 5413 4697 5451 4731
rect 5485 4697 5523 4731
rect 5557 4697 5595 4731
rect 5629 4697 5667 4731
rect 5701 4697 5739 4731
rect 5773 4697 5811 4731
rect 5845 4697 5883 4731
rect 5917 4697 5955 4731
rect 5989 4697 6027 4731
rect 6061 4697 6099 4731
rect 6133 4697 6171 4731
rect 6205 4697 6243 4731
rect 6277 4697 6315 4731
rect 6349 4697 6387 4731
rect 6421 4697 6459 4731
rect 6493 4697 6531 4731
rect 6565 4697 6603 4731
rect 6637 4697 6675 4731
rect 6709 4697 6747 4731
rect 6781 4697 6819 4731
rect 6853 4697 6891 4731
rect 6925 4697 6963 4731
rect 6997 4697 7035 4731
rect 7069 4697 7107 4731
rect 7141 4697 7179 4731
rect 7213 4697 7251 4731
rect 7285 4697 7323 4731
rect 7357 4697 7395 4731
rect 7429 4697 7467 4731
rect 7501 4697 7539 4731
rect 7573 4697 7611 4731
rect 7645 4697 7683 4731
rect 7717 4697 7755 4731
rect 7789 4697 7827 4731
rect 7861 4697 7899 4731
rect 7933 4697 7971 4731
rect 8005 4697 8043 4731
rect 3366 4659 8043 4697
rect 3366 4625 3444 4659
rect 3478 4625 3517 4659
rect 3551 4625 3590 4659
rect 3624 4625 3663 4659
rect 3697 4625 3736 4659
rect 3770 4625 3809 4659
rect 3843 4625 3882 4659
rect 3916 4625 3955 4659
rect 3989 4625 4028 4659
rect 4062 4625 4101 4659
rect 4135 4625 4174 4659
rect 4208 4625 4247 4659
rect 4281 4625 4320 4659
rect 4354 4625 4393 4659
rect 4427 4625 4466 4659
rect 4500 4625 4539 4659
rect 4573 4625 4612 4659
rect 4646 4625 4685 4659
rect 4719 4625 4758 4659
rect 4792 4625 4831 4659
rect 4865 4625 4904 4659
rect 4938 4625 4977 4659
rect 5011 4625 5050 4659
rect 5084 4625 5123 4659
rect 5157 4625 5196 4659
rect 5230 4625 5269 4659
rect 5303 4625 5342 4659
rect 5376 4625 5415 4659
rect 5449 4625 5488 4659
rect 5522 4625 5561 4659
rect 5595 4625 5634 4659
rect 5668 4625 5707 4659
rect 5741 4625 5780 4659
rect 5814 4625 5853 4659
rect 5887 4625 5926 4659
rect 5960 4625 5999 4659
rect 6033 4625 6072 4659
rect 6106 4625 6145 4659
rect 6179 4625 6218 4659
rect 6252 4625 6291 4659
rect 6325 4625 6364 4659
rect 6398 4625 6437 4659
rect 6471 4625 6510 4659
rect 6544 4625 6583 4659
rect 6617 4625 6656 4659
rect 6690 4625 6729 4659
rect 6763 4625 6802 4659
rect 6836 4625 6875 4659
rect 6909 4625 6948 4659
rect 6982 4625 7021 4659
rect 7055 4625 7094 4659
rect 7128 4625 7167 4659
rect 7201 4625 7240 4659
rect 7274 4625 7313 4659
rect 7347 4625 7386 4659
rect 7420 4625 7459 4659
rect 7493 4625 7532 4659
rect 7566 4625 7605 4659
rect 7639 4625 7678 4659
rect 7712 4625 7751 4659
rect 7785 4625 7824 4659
rect 7858 4625 7897 4659
rect 7931 4625 7970 4659
rect 8004 4625 8043 4659
rect 13333 4625 13367 4731
rect 3366 4619 13367 4625
rect 3366 4613 3484 4619
rect 3366 4579 3372 4613
rect 3406 4582 3484 4613
tri 3484 4594 3509 4619 nw
rect 3406 4579 3444 4582
rect 3366 4548 3444 4579
rect 3478 4548 3484 4582
rect 3366 4537 3484 4548
rect 3366 4503 3372 4537
rect 3406 4505 3484 4537
rect 3406 4503 3444 4505
rect 3366 4471 3444 4503
rect 3478 4471 3484 4505
rect 3366 4461 3484 4471
rect 3366 4427 3372 4461
rect 3406 4428 3484 4461
rect 3406 4427 3444 4428
rect 3366 4394 3444 4427
rect 3478 4394 3484 4428
rect 3366 4384 3484 4394
rect 3366 4350 3372 4384
rect 3406 4351 3484 4384
rect 3406 4350 3444 4351
rect 3366 4317 3444 4350
rect 3478 4317 3484 4351
rect 3366 4307 3484 4317
rect 3366 4273 3372 4307
rect 3406 4274 3484 4307
rect 6930 4283 13084 4463
rect 3406 4273 3444 4274
rect 3366 4240 3444 4273
rect 3478 4240 3484 4274
rect 3366 4230 3484 4240
rect 3366 4196 3372 4230
rect 3406 4197 3484 4230
rect 3406 4196 3444 4197
rect 3366 4163 3444 4196
rect 3478 4163 3484 4197
rect 3366 4153 3484 4163
rect 3366 4119 3372 4153
rect 3406 4120 3484 4153
rect 3406 4119 3444 4120
rect 3366 4086 3444 4119
rect 3478 4086 3484 4120
rect 3366 4076 3484 4086
rect 3366 4042 3372 4076
rect 3406 4043 3484 4076
rect 16105 4176 16877 4188
rect 16105 4142 16111 4176
rect 16145 4142 16287 4176
rect 16321 4142 16463 4176
rect 16497 4142 16639 4176
rect 16673 4142 16837 4176
rect 16871 4142 16877 4176
rect 16105 4104 16877 4142
rect 16105 4070 16111 4104
rect 16145 4070 16287 4104
rect 16321 4070 16463 4104
rect 16497 4070 16639 4104
rect 16673 4070 16837 4104
rect 16871 4070 16877 4104
rect 16105 4058 16877 4070
rect 3406 4042 3444 4043
rect 3366 4009 3444 4042
rect 3478 4009 3484 4043
tri 17329 4030 17354 4055 se
rect 17354 4030 17552 4234
tri 17552 4209 17577 4234 nw
tri 17633 4209 17658 4234 ne
tri 17552 4030 17577 4055 sw
tri 17633 4030 17658 4055 se
rect 17658 4030 17856 4234
tri 17856 4209 17881 4234 nw
tri 17928 4209 17953 4234 ne
tri 17856 4030 17881 4055 sw
tri 17928 4030 17953 4055 se
rect 17953 4030 18151 4234
tri 18151 4209 18176 4234 nw
tri 18151 4030 18176 4055 sw
rect 3366 3999 3484 4009
rect 3366 3965 3372 3999
rect 3406 3966 3484 3999
rect 3406 3965 3444 3966
tri 3345 3932 3366 3953 se
rect 3366 3932 3444 3965
rect 3478 3932 3484 3966
tri 3341 3928 3345 3932 se
rect 3345 3928 3484 3932
rect 23 3922 3484 3928
rect 23 3888 35 3922
rect 69 3888 108 3922
rect 142 3888 181 3922
rect 215 3888 254 3922
rect 288 3888 327 3922
rect 361 3888 400 3922
rect 434 3888 473 3922
rect 507 3888 546 3922
rect 580 3888 619 3922
rect 653 3888 692 3922
rect 726 3888 765 3922
rect 799 3888 838 3922
rect 872 3888 911 3922
rect 945 3888 984 3922
rect 1018 3888 1057 3922
rect 1091 3888 1130 3922
rect 1164 3888 1203 3922
rect 1237 3888 1276 3922
rect 1310 3888 1349 3922
rect 1383 3888 1422 3922
rect 1456 3888 1495 3922
rect 1529 3888 1568 3922
rect 1602 3888 1641 3922
rect 1675 3888 1714 3922
rect 1748 3888 1787 3922
rect 1821 3888 1860 3922
rect 1894 3888 1932 3922
rect 1966 3888 2004 3922
rect 2038 3888 2076 3922
rect 2110 3888 2148 3922
rect 2182 3888 2220 3922
rect 2254 3888 2292 3922
rect 2326 3888 2364 3922
rect 2398 3888 2436 3922
rect 2470 3888 2508 3922
rect 2542 3888 2580 3922
rect 2614 3888 2652 3922
rect 2686 3888 2724 3922
rect 2758 3888 2796 3922
rect 2830 3888 2868 3922
rect 2902 3888 2940 3922
rect 2974 3888 3012 3922
rect 3046 3888 3084 3922
rect 3118 3888 3156 3922
rect 3190 3888 3228 3922
rect 3262 3888 3300 3922
rect 3334 3888 3372 3922
rect 3406 3888 3484 3922
rect 23 3854 3444 3888
rect 3478 3854 3484 3888
rect 23 3850 3484 3854
rect 23 3816 35 3850
rect 69 3816 109 3850
rect 143 3816 183 3850
rect 217 3816 257 3850
rect 291 3816 331 3850
rect 365 3816 405 3850
rect 439 3816 479 3850
rect 513 3816 553 3850
rect 587 3816 627 3850
rect 661 3816 701 3850
rect 735 3816 775 3850
rect 809 3816 849 3850
rect 883 3816 923 3850
rect 957 3816 996 3850
rect 1030 3816 1069 3850
rect 1103 3816 1142 3850
rect 1176 3816 1215 3850
rect 1249 3816 1288 3850
rect 1322 3816 1361 3850
rect 1395 3816 1434 3850
rect 1468 3816 1507 3850
rect 1541 3816 1580 3850
rect 1614 3816 1653 3850
rect 1687 3816 1726 3850
rect 1760 3816 1799 3850
rect 1833 3816 1872 3850
rect 1906 3816 1945 3850
rect 1979 3816 2018 3850
rect 2052 3816 2091 3850
rect 2125 3816 2164 3850
rect 2198 3816 2237 3850
rect 2271 3816 2310 3850
rect 2344 3816 2383 3850
rect 2417 3816 2456 3850
rect 2490 3816 2529 3850
rect 2563 3816 2602 3850
rect 2636 3816 2675 3850
rect 2709 3816 2748 3850
rect 2782 3816 2821 3850
rect 2855 3816 2894 3850
rect 2928 3816 2967 3850
rect 3001 3816 3040 3850
rect 3074 3816 3113 3850
rect 3147 3816 3186 3850
rect 3220 3816 3259 3850
rect 3293 3816 3332 3850
rect 3366 3816 3484 3850
rect 23 3810 3484 3816
rect 13494 3774 13500 3954
rect 13680 3838 13686 3954
rect 13616 3774 13622 3838
rect 15793 3754 17001 4030
tri 13232 3720 13238 3726 se
rect 13238 3720 15927 3726
rect 15929 3725 15957 3726
tri 13198 3686 13232 3720 se
rect 13232 3686 15927 3720
tri 13196 3684 13198 3686 se
rect 13198 3684 15927 3686
tri 13158 3646 13196 3684 se
rect 13196 3646 15927 3684
tri 13124 3612 13158 3646 se
rect 13158 3612 15927 3646
tri 13054 3542 13124 3612 se
rect 13124 3606 15927 3612
rect 15928 3607 15958 3725
rect 15959 3720 16597 3726
rect 15959 3686 16199 3720
rect 16233 3686 16551 3720
rect 16585 3686 16597 3720
rect 15929 3606 15957 3607
rect 15959 3606 16597 3686
rect 16912 3718 16970 3724
rect 16912 3684 16924 3718
rect 16958 3684 16970 3718
rect 16912 3646 16970 3684
rect 16912 3612 16924 3646
rect 16958 3638 16970 3646
tri 16970 3638 16995 3663 sw
rect 16958 3612 17189 3638
rect 16912 3606 17189 3612
rect 13124 3542 13238 3606
tri 13238 3542 13302 3606 nw
tri 12986 3474 13054 3542 se
rect 13054 3474 13170 3542
tri 13170 3474 13238 3542 nw
rect 18093 3532 18479 3578
rect 6446 3459 13039 3474
rect 6446 3343 6452 3459
rect 6568 3343 13039 3459
tri 13039 3343 13170 3474 nw
rect 13789 3427 14333 3504
rect 13789 3375 13882 3427
rect 13934 3375 14333 3427
rect 13789 3363 14333 3375
rect 10314 3197 12997 3315
rect 13789 3311 13818 3363
rect 13870 3311 13882 3363
rect 13934 3311 14333 3363
rect 13789 3263 14333 3311
rect 10314 3137 12937 3197
tri 12937 3137 12997 3197 nw
rect 13112 3147 13432 3153
rect 10314 3103 12903 3137
tri 12903 3103 12937 3137 nw
rect 10314 3099 12899 3103
tri 12899 3099 12903 3103 nw
rect 10314 3039 12882 3099
tri 12882 3082 12899 3099 nw
rect 13164 3143 13432 3147
tri 13432 3143 13442 3153 sw
rect 13164 3137 19133 3143
rect 13164 3125 13425 3137
rect 13164 3103 13167 3125
tri 13167 3103 13189 3125 nw
tri 13385 3103 13407 3125 ne
rect 13407 3103 13425 3125
rect 13459 3103 13498 3137
rect 13532 3103 13571 3137
rect 13605 3103 13644 3137
rect 13678 3103 13717 3137
rect 13751 3103 13790 3137
rect 13824 3103 13863 3137
rect 13897 3103 13936 3137
rect 13970 3103 14009 3137
rect 14043 3103 14082 3137
rect 14116 3103 14155 3137
rect 14189 3103 14228 3137
rect 14262 3103 14301 3137
rect 14335 3103 14374 3137
rect 14408 3103 14447 3137
rect 14481 3103 14519 3137
rect 14553 3103 14591 3137
rect 14625 3103 14663 3137
rect 14697 3103 14735 3137
rect 14769 3103 14807 3137
rect 14841 3103 14879 3137
rect 14913 3103 14951 3137
rect 14985 3103 15023 3137
rect 15057 3103 15095 3137
rect 15129 3103 15167 3137
rect 15201 3103 15239 3137
rect 15273 3103 15311 3137
rect 15345 3103 15383 3137
rect 15417 3103 15455 3137
rect 15489 3103 15527 3137
rect 15561 3103 15599 3137
rect 15633 3103 15671 3137
rect 15705 3103 15743 3137
rect 15777 3103 15815 3137
rect 15849 3103 15887 3137
rect 15921 3103 15959 3137
rect 15993 3103 16031 3137
rect 16065 3103 16103 3137
rect 16137 3103 16175 3137
rect 16209 3103 16247 3137
rect 16281 3103 16319 3137
rect 16353 3103 16391 3137
rect 16425 3103 16463 3137
rect 16497 3103 16535 3137
rect 16569 3103 16607 3137
rect 16641 3103 16679 3137
rect 16713 3103 16751 3137
rect 16785 3103 16823 3137
rect 16857 3103 16895 3137
rect 16929 3103 16967 3137
rect 17001 3103 17039 3137
rect 17073 3103 17111 3137
rect 17145 3103 17183 3137
rect 17217 3103 17255 3137
rect 17289 3103 17327 3137
rect 17361 3103 17399 3137
rect 17433 3103 17471 3137
rect 17505 3103 17543 3137
rect 17577 3103 17615 3137
rect 17649 3103 17687 3137
rect 17721 3103 17759 3137
rect 17793 3103 17831 3137
rect 17865 3103 17903 3137
rect 17937 3103 17975 3137
rect 18009 3103 18047 3137
rect 18081 3103 18119 3137
rect 18153 3103 18191 3137
rect 18225 3103 18263 3137
rect 18297 3103 18335 3137
rect 18369 3103 18407 3137
rect 18441 3103 18479 3137
rect 18513 3103 18551 3137
rect 18585 3103 18623 3137
rect 18657 3103 18695 3137
rect 18729 3103 18767 3137
rect 18801 3103 18839 3137
rect 18873 3103 18911 3137
rect 18945 3103 18983 3137
rect 19017 3103 19133 3137
tri 13164 3100 13167 3103 nw
tri 13407 3100 13410 3103 ne
rect 13410 3100 19133 3103
tri 13410 3099 13411 3100 ne
rect 13411 3099 19133 3100
tri 13411 3097 13413 3099 ne
rect 13413 3097 19093 3099
rect 13112 3083 13164 3095
rect 10314 3023 11009 3039
tri 11009 3023 11025 3039 nw
tri 12740 3023 12756 3039 ne
rect 12756 3023 12882 3039
rect 13210 3045 13216 3097
rect 13268 3045 13280 3097
rect 13332 3069 13338 3097
tri 13338 3069 13366 3097 sw
tri 19051 3069 19079 3097 ne
rect 19079 3069 19093 3097
rect 13332 3065 18278 3069
tri 18278 3065 18282 3069 sw
tri 19079 3065 19083 3069 ne
rect 19083 3065 19093 3069
rect 19127 3065 19133 3099
rect 13332 3064 18282 3065
tri 18282 3064 18283 3065 sw
tri 19083 3064 19084 3065 ne
rect 19084 3064 19133 3065
rect 13332 3045 18283 3064
rect 13210 3041 18283 3045
rect 13112 3025 13164 3031
tri 18265 3025 18281 3041 ne
rect 18281 3025 18283 3041
tri 18281 3023 18283 3025 ne
tri 18283 3023 18324 3064 sw
tri 19084 3061 19087 3064 ne
rect 19087 3023 19133 3064
rect 10314 2989 10975 3023
tri 10975 2989 11009 3023 nw
tri 12756 2989 12790 3023 ne
rect 12790 2989 12882 3023
tri 18283 3013 18293 3023 ne
rect 18293 3013 18324 3023
rect 10314 2947 10933 2989
tri 10933 2947 10975 2989 nw
tri 12790 2947 12832 2989 ne
rect 12832 2947 12882 2989
rect 10314 2913 10899 2947
tri 10899 2913 10933 2947 nw
tri 12832 2913 12866 2947 ne
rect 12866 2913 12882 2947
rect 10314 2872 10858 2913
tri 10858 2872 10899 2913 nw
tri 12866 2897 12882 2913 ne
rect 13286 3008 18251 3013
tri 18251 3008 18256 3013 sw
tri 18293 3008 18298 3013 ne
rect 18298 3008 18324 3013
rect 13286 3007 18256 3008
rect 13338 2989 18256 3007
tri 18256 2989 18275 3008 sw
tri 18298 2989 18317 3008 ne
rect 18317 2989 18324 3008
tri 18324 2989 18358 3023 sw
rect 19087 2989 19093 3023
rect 19127 2989 19133 3023
rect 13338 2985 18275 2989
tri 13338 2960 13363 2985 nw
tri 18238 2967 18256 2985 ne
rect 18256 2982 18275 2985
tri 18275 2982 18282 2989 sw
tri 18317 2982 18324 2989 ne
rect 18324 2982 18358 2989
tri 18358 2982 18365 2989 sw
rect 18256 2967 18282 2982
tri 18282 2967 18297 2982 sw
tri 18324 2967 18339 2982 ne
rect 18339 2967 18956 2982
tri 18256 2960 18263 2967 ne
rect 18263 2960 18297 2967
rect 13286 2943 13338 2955
tri 18263 2947 18276 2960 ne
rect 18276 2954 18297 2960
tri 18297 2954 18310 2967 sw
tri 18339 2954 18352 2967 ne
rect 18352 2962 18956 2967
tri 18956 2962 18976 2982 sw
rect 18352 2954 18976 2962
rect 18276 2947 18310 2954
tri 18310 2947 18317 2954 sw
tri 18943 2947 18950 2954 ne
rect 18950 2947 18976 2954
tri 18976 2947 18991 2962 sw
rect 19087 2947 19133 2989
tri 18276 2926 18297 2947 ne
rect 18297 2926 18317 2947
tri 18317 2926 18338 2947 sw
tri 18950 2926 18971 2947 ne
rect 18971 2926 18991 2947
tri 18297 2913 18310 2926 ne
rect 18310 2925 18910 2926
tri 18910 2925 18911 2926 sw
tri 18971 2925 18972 2926 ne
rect 18972 2925 18991 2926
rect 18310 2921 18911 2925
tri 18911 2921 18915 2925 sw
tri 18972 2921 18976 2925 ne
rect 18976 2921 18991 2925
tri 18991 2921 19017 2947 sw
rect 18310 2913 18915 2921
tri 18915 2913 18923 2921 sw
tri 18976 2913 18984 2921 ne
rect 18984 2913 19017 2921
tri 18310 2898 18325 2913 ne
rect 18325 2898 18923 2913
rect 13286 2885 13338 2891
tri 18897 2885 18910 2898 ne
rect 18910 2885 18923 2898
tri 18910 2884 18911 2885 ne
rect 18911 2884 18923 2885
tri 18923 2884 18952 2913 sw
tri 18984 2908 18989 2913 ne
tri 18911 2872 18923 2884 ne
rect 18923 2872 18952 2884
rect 10314 2838 10824 2872
tri 10824 2838 10858 2872 nw
tri 18923 2871 18924 2872 ne
rect 10314 2797 10783 2838
tri 10783 2797 10824 2838 nw
rect 10314 2763 10749 2797
tri 10749 2763 10783 2797 nw
rect 10314 2722 10708 2763
tri 10708 2722 10749 2763 nw
rect 12956 2736 12962 2852
rect 13078 2838 13084 2852
tri 13084 2838 13098 2852 sw
rect 13078 2797 13098 2838
tri 13098 2797 13139 2838 sw
rect 13078 2789 13139 2797
tri 13139 2789 13147 2797 sw
rect 13078 2763 15337 2789
tri 15337 2763 15363 2789 sw
rect 13078 2745 15363 2763
tri 15363 2745 15381 2763 sw
rect 13078 2736 15381 2745
tri 15298 2722 15312 2736 ne
rect 15312 2722 15381 2736
rect 10314 2688 10674 2722
tri 10674 2688 10708 2722 nw
tri 15312 2711 15323 2722 ne
rect 15323 2707 15381 2722
rect 18924 2702 18952 2872
rect 18989 2702 19017 2913
rect 19087 2913 19093 2947
rect 19127 2913 19133 2947
rect 19087 2872 19133 2913
rect 19087 2838 19093 2872
rect 19127 2838 19133 2872
rect 19087 2797 19133 2838
rect 19087 2763 19093 2797
rect 19127 2763 19133 2797
rect 19087 2722 19133 2763
rect 10314 2647 10633 2688
tri 10633 2647 10674 2688 nw
rect 10314 2613 10599 2647
tri 10599 2613 10633 2647 nw
tri 12714 2613 12742 2641 se
rect 10314 2400 10590 2613
tri 10590 2604 10599 2613 nw
tri 12705 2604 12714 2613 se
rect 12714 2604 12742 2613
tri 12673 2572 12705 2604 se
rect 12705 2584 12742 2604
rect 12705 2572 12882 2584
rect 13366 2580 13372 2696
rect 13488 2688 14358 2696
tri 14358 2688 14366 2696 sw
rect 19087 2688 19093 2722
rect 19127 2688 19133 2722
rect 13488 2647 14366 2688
tri 14366 2647 14407 2688 sw
rect 19087 2647 19133 2688
rect 13488 2645 14407 2647
tri 14407 2645 14409 2647 sw
rect 13488 2580 14409 2645
tri 14254 2572 14262 2580 ne
rect 14262 2572 14409 2580
tri 12646 2545 12673 2572 se
rect 12673 2545 12882 2572
tri 14262 2555 14279 2572 ne
rect 14279 2534 14409 2572
rect 17108 2621 17160 2627
rect 17108 2557 17160 2569
rect 17108 2499 17160 2505
tri 17108 2497 17110 2499 ne
rect 17110 2497 17160 2499
tri 17110 2493 17114 2497 ne
rect 17114 2493 17160 2497
rect 19087 2613 19093 2647
rect 19127 2613 19133 2647
rect 19087 2572 19133 2613
rect 19087 2538 19093 2572
rect 19127 2538 19133 2572
rect 19087 2497 19133 2538
rect 19087 2463 19093 2497
rect 19127 2463 19133 2497
rect 19087 2451 19133 2463
rect 10314 2183 10432 2400
tri 10432 2340 10492 2400 nw
tri 10432 2183 10492 2243 sw
rect 10691 2234 10697 2350
rect 10877 2234 10883 2350
rect 10314 1580 10590 2183
rect 12882 2086 13072 2286
rect 18988 2271 19106 2283
rect 11578 1872 11838 2050
tri 11578 1870 11580 1872 ne
rect 11580 1870 11836 1872
tri 11836 1870 11838 1872 nw
tri 17108 1812 17114 1818 se
rect 17114 1812 17160 1818
rect 17108 1806 17160 1812
rect 17108 1742 17160 1754
tri 10590 1580 10732 1722 sw
rect 17108 1684 17160 1690
tri 17108 1678 17114 1684 ne
rect 17114 1678 17160 1684
rect 13286 1617 13338 1623
rect 10314 1488 10432 1580
tri 10432 1488 10524 1580 nw
tri 13261 1547 13286 1572 se
rect 13286 1553 13338 1565
rect 10835 1495 10841 1547
rect 10893 1495 10905 1547
rect 10957 1501 13286 1547
rect 10957 1495 13338 1501
rect 10613 1426 13164 1432
rect 10613 1392 10657 1426
rect 10691 1392 10730 1426
rect 10764 1392 10803 1426
rect 10837 1392 10876 1426
rect 10910 1392 10949 1426
rect 10983 1392 11022 1426
rect 11056 1392 11095 1426
rect 11129 1392 11168 1426
rect 11202 1392 11241 1426
rect 11275 1392 11314 1426
rect 11348 1392 11387 1426
rect 11421 1392 11460 1426
rect 11494 1392 11533 1426
rect 11567 1392 11606 1426
rect 11640 1392 11678 1426
rect 11712 1392 11750 1426
rect 11784 1392 11822 1426
rect 11856 1392 11894 1426
rect 11928 1392 11966 1426
rect 12000 1392 12038 1426
rect 12072 1392 12110 1426
rect 12144 1392 12182 1426
rect 12216 1392 12254 1426
rect 12288 1392 12326 1426
rect 12360 1392 12398 1426
rect 12432 1392 12470 1426
rect 12504 1392 12542 1426
rect 12576 1392 12614 1426
rect 12648 1392 12686 1426
rect 12720 1392 12758 1426
rect 12792 1392 12830 1426
rect 12864 1392 12902 1426
rect 12936 1392 12974 1426
rect 13008 1392 13046 1426
rect 13080 1392 13112 1426
rect 10613 1386 13112 1392
rect 10613 1328 10953 1386
tri 10953 1333 11006 1386 nw
tri 13087 1361 13112 1386 ne
rect 13112 1362 13164 1374
rect 10613 1322 10807 1328
rect 10613 1316 10691 1322
rect 10613 1282 10619 1316
rect 10653 1282 10691 1316
rect 10613 1244 10691 1282
rect 10613 1210 10619 1244
rect 10653 1210 10691 1244
rect 10613 1172 10691 1210
rect 10613 1138 10619 1172
rect 10653 1142 10691 1172
rect 13112 1304 13164 1310
rect 10653 1138 10807 1142
rect 18988 1301 18994 2271
rect 19100 1301 19106 2271
rect 18988 1262 19106 1301
rect 18988 1228 18994 1262
rect 19028 1228 19066 1262
rect 19100 1228 19106 1262
rect 18988 1189 19106 1228
rect 18988 1155 18994 1189
rect 19028 1155 19066 1189
rect 19100 1155 19106 1189
rect 10613 1136 10807 1138
rect 10613 1100 10691 1136
rect 10613 1066 10619 1100
rect 10653 1066 10691 1100
rect 13442 1089 13448 1141
rect 13500 1089 13506 1141
rect 18988 1116 19106 1155
rect 10613 1028 10691 1066
rect 10613 994 10619 1028
rect 10653 994 10691 1028
rect 18988 1082 18994 1116
rect 19028 1082 19066 1116
rect 19100 1082 19106 1116
rect 18988 1043 19106 1082
rect 18988 1009 18994 1043
rect 19028 1009 19066 1043
rect 19100 1009 19106 1043
rect 10613 956 10691 994
rect 10613 922 10619 956
rect 10653 922 10691 956
rect 10613 884 10691 922
tri 10953 982 10978 1007 sw
tri 13153 982 13171 1000 se
rect 13171 982 13262 1000
rect 10953 936 11523 982
rect 11824 942 13262 982
rect 13442 945 13448 997
rect 13500 945 13506 997
rect 18988 970 19106 1009
rect 11824 936 13173 942
tri 13173 936 13179 942 nw
rect 18988 936 18994 970
rect 19028 936 19066 970
rect 19100 936 19106 970
tri 10953 911 10978 936 nw
rect 18988 924 19106 936
rect 10613 850 10619 884
rect 10653 850 10691 884
rect 10613 812 10691 850
rect 10613 778 10619 812
rect 10653 778 10691 812
rect 10613 740 10691 778
rect 10613 706 10619 740
rect 10653 706 10691 740
tri 18937 833 18988 884 se
rect 18988 833 19009 924
rect 10613 668 10691 706
rect 10613 634 10619 668
rect 10653 634 10691 668
rect 13442 657 13448 709
rect 13500 657 13506 709
tri 17108 673 17114 679 se
rect 17114 673 17160 679
rect 17108 667 17160 673
rect 10613 596 10691 634
rect 10613 562 10619 596
rect 10653 562 10691 596
rect 15111 611 15163 617
rect 10613 524 10691 562
tri 12458 550 12476 568 se
rect 12476 550 13262 568
rect 10613 490 10619 524
rect 10653 490 10691 524
rect 11824 510 13262 550
rect 13442 513 13448 565
rect 13500 513 13506 565
rect 15111 547 15163 559
rect 11824 504 12478 510
tri 12478 504 12484 510 nw
rect 10613 452 10691 490
rect 10613 418 10619 452
rect 10653 418 10691 452
rect 11523 494 11566 504
tri 11566 494 11576 504 nw
rect 17108 603 17160 615
rect 17108 545 17160 551
rect 10613 380 10691 418
tri 11503 413 11523 433 se
rect 11523 413 11551 494
tri 11551 479 11566 494 nw
rect 15111 489 15163 495
tri 18184 479 18185 480 ne
rect 18185 479 18460 480
tri 18185 460 18204 479 ne
rect 18204 460 18460 479
tri 18204 438 18226 460 ne
rect 18226 438 18460 460
tri 11551 413 11576 438 sw
tri 18226 413 18251 438 ne
rect 18251 413 18460 438
tri 11498 408 11503 413 se
rect 11503 408 11551 413
tri 18251 408 18256 413 ne
rect 18256 408 18460 413
tri 18256 402 18262 408 ne
rect 10613 346 10619 380
rect 10653 346 10691 380
rect 18262 379 18460 408
tri 18460 379 18461 380 sw
tri 18936 379 18937 380 se
rect 18937 379 19009 833
tri 19009 827 19106 924 nw
rect 19108 737 19154 749
rect 19108 703 19114 737
rect 19148 703 19154 737
rect 19108 656 19154 703
rect 19108 622 19114 656
rect 19148 622 19154 656
rect 19108 575 19154 622
rect 19108 541 19114 575
rect 19148 541 19154 575
rect 19108 494 19154 541
rect 10613 332 10691 346
tri 10691 332 10735 376 sw
rect 18262 355 18461 379
tri 18461 355 18485 379 sw
tri 18912 355 18936 379 se
rect 18936 355 19009 379
rect 10613 308 10735 332
rect 10613 274 10619 308
rect 10653 298 10735 308
tri 10735 298 10769 332 sw
rect 18262 316 19009 355
tri 19033 298 19048 313 se
rect 19048 298 19080 480
rect 10653 274 10769 298
rect 10613 251 10769 274
tri 10769 251 10816 298 sw
tri 19023 288 19033 298 se
rect 19033 288 19080 298
rect 10613 236 10816 251
tri 10816 236 10831 251 sw
rect 18101 236 18107 288
rect 18159 236 18171 288
rect 18223 274 19080 288
rect 18223 251 19057 274
tri 19057 251 19080 274 nw
rect 19108 460 19114 494
rect 19148 460 19154 494
rect 19108 413 19154 460
rect 19108 379 19114 413
rect 19148 379 19154 413
rect 19108 332 19154 379
rect 19108 298 19114 332
rect 19148 298 19154 332
rect 19108 251 19154 298
rect 18223 236 19042 251
tri 19042 236 19057 251 nw
rect 10613 235 17934 236
rect 10613 201 10619 235
rect 10653 208 17934 235
rect 10653 201 13824 208
rect 10613 162 13824 201
rect 10613 128 10619 162
rect 10653 156 13824 162
rect 13876 156 13917 208
rect 13969 156 14010 208
rect 14062 207 17214 208
rect 14062 156 15117 207
rect 10653 155 15117 156
rect 15169 155 17214 207
rect 10653 144 17214 155
rect 10653 128 13824 144
rect 10613 124 13824 128
rect 13876 124 13917 144
rect 13969 124 14010 144
rect 14062 143 17214 144
rect 14062 124 15117 143
rect 15169 124 17214 143
rect 17330 130 17934 208
rect 19108 217 19114 251
rect 19148 217 19154 251
tri 17934 130 17978 174 sw
rect 19108 130 19154 217
rect 17330 124 19154 130
rect 10613 90 10729 124
rect 10763 90 10801 124
rect 10835 90 10873 124
rect 10907 90 10945 124
rect 10979 90 11017 124
rect 11051 90 11089 124
rect 11123 90 11161 124
rect 11195 90 11233 124
rect 11267 90 11305 124
rect 11339 90 11377 124
rect 11411 90 11449 124
rect 11483 90 11521 124
rect 11555 90 11593 124
rect 11627 90 11665 124
rect 11699 90 11737 124
rect 11771 90 11809 124
rect 11843 90 11881 124
rect 11915 90 11953 124
rect 11987 90 12025 124
rect 12059 90 12097 124
rect 12131 90 12169 124
rect 12203 90 12241 124
rect 12275 90 12313 124
rect 12347 90 12385 124
rect 12419 90 12457 124
rect 12491 90 12529 124
rect 12563 90 12601 124
rect 12635 90 12673 124
rect 12707 90 12745 124
rect 12779 90 12817 124
rect 12851 90 12889 124
rect 12923 90 12961 124
rect 12995 90 13033 124
rect 13067 90 13105 124
rect 13139 90 13177 124
rect 13211 90 13249 124
rect 13283 90 13321 124
rect 13355 90 13393 124
rect 13427 90 13465 124
rect 13499 90 13537 124
rect 13571 90 13609 124
rect 13643 90 13681 124
rect 13715 90 13753 124
rect 13787 92 13824 124
rect 13876 92 13897 124
rect 13787 90 13825 92
rect 13859 90 13897 92
rect 13931 90 13969 92
rect 14003 92 14010 124
rect 14003 90 14041 92
rect 14075 90 14113 124
rect 14147 90 14185 124
rect 14219 90 14258 124
rect 14292 90 14331 124
rect 14365 90 14404 124
rect 14438 90 14477 124
rect 14511 90 14550 124
rect 14584 90 14623 124
rect 14657 90 14696 124
rect 14730 90 14769 124
rect 14803 90 14842 124
rect 14876 90 14915 124
rect 14949 90 14988 124
rect 15022 90 15061 124
rect 15095 91 15117 124
rect 15169 91 15207 124
rect 15095 90 15134 91
rect 15168 90 15207 91
rect 15241 90 15280 124
rect 15314 90 15353 124
rect 15387 90 15426 124
rect 15460 90 15499 124
rect 15533 90 15572 124
rect 15606 90 15645 124
rect 15679 90 15718 124
rect 15752 90 15791 124
rect 15825 90 15864 124
rect 15898 90 15937 124
rect 15971 90 16010 124
rect 16044 90 16083 124
rect 16117 90 16156 124
rect 16190 90 16229 124
rect 16263 90 16302 124
rect 16336 90 16375 124
rect 16409 90 16448 124
rect 16482 90 16521 124
rect 16555 90 16594 124
rect 16628 90 16667 124
rect 16701 90 16740 124
rect 16774 90 16813 124
rect 16847 90 16886 124
rect 16920 90 16959 124
rect 16993 90 17032 124
rect 17066 90 17105 124
rect 17139 90 17178 124
rect 17212 92 17214 124
rect 17212 90 17251 92
rect 17285 90 17324 92
rect 17358 90 17397 124
rect 17431 90 17470 124
rect 17504 90 17543 124
rect 17577 90 17616 124
rect 17650 90 17689 124
rect 17723 90 17762 124
rect 17796 90 17835 124
rect 17869 90 17908 124
rect 17942 90 17981 124
rect 18015 90 18054 124
rect 18088 90 18127 124
rect 18161 90 18200 124
rect 18234 90 18273 124
rect 18307 90 18346 124
rect 18380 90 18419 124
rect 18453 90 18492 124
rect 18526 90 18565 124
rect 18599 90 18638 124
rect 18672 90 18711 124
rect 18745 90 18784 124
rect 18818 90 18857 124
rect 18891 90 18930 124
rect 18964 90 19003 124
rect 19037 90 19076 124
rect 19110 90 19154 124
rect 10613 84 19154 90
<< rmetal1 >>
rect 6560 6416 6562 6417
rect 6560 6302 6561 6416
rect 6560 6301 6562 6302
rect 6598 6416 6600 6417
rect 6599 6302 6600 6416
rect 6598 6301 6600 6302
rect 6846 6337 6892 6338
rect 6846 6336 6847 6337
rect 6891 6336 6892 6337
rect 6846 6299 6847 6300
rect 6891 6299 6892 6300
rect 6846 6298 6892 6299
rect 6846 6080 6892 6081
rect 6846 6079 6847 6080
rect 6891 6079 6892 6080
rect 6846 6042 6847 6043
rect 6891 6042 6892 6043
rect 6846 6041 6892 6042
rect 6846 5644 6892 5645
rect 6846 5643 6847 5644
rect 6891 5643 6892 5644
rect 6846 5612 6847 5613
rect 6891 5612 6892 5613
rect 6846 5611 6892 5612
rect 6846 5308 6892 5309
rect 6846 5307 6847 5308
rect 6891 5307 6892 5308
rect 6846 5276 6847 5277
rect 6891 5276 6892 5277
rect 6846 5275 6892 5276
rect 9856 6172 9858 6173
rect 9894 6172 9896 6173
rect 9856 6128 9857 6172
rect 9895 6128 9896 6172
rect 9856 6127 9858 6128
rect 9894 6127 9896 6128
rect 9856 5824 9858 5825
rect 9894 5824 9896 5825
rect 9856 5780 9857 5824
rect 9895 5780 9896 5824
rect 9856 5779 9858 5780
rect 9894 5779 9896 5780
rect 9856 5476 9858 5477
rect 9894 5476 9896 5477
rect 9856 5432 9857 5476
rect 9895 5432 9896 5476
rect 9856 5431 9858 5432
rect 9894 5431 9896 5432
rect 6780 5171 6782 5172
rect 6780 5127 6781 5171
rect 6780 5126 6782 5127
rect 6812 5171 6814 5172
rect 6813 5127 6814 5171
rect 6812 5126 6814 5127
rect 6920 5084 9833 5085
rect 6920 5083 6921 5084
rect 9832 5083 9833 5084
rect 6920 5054 6921 5055
rect 9832 5054 9833 5055
rect 6920 5053 9833 5054
rect 10115 6172 10117 6173
rect 10153 6172 10155 6173
rect 10115 6128 10116 6172
rect 10154 6128 10155 6172
rect 10115 6127 10117 6128
rect 10153 6127 10155 6128
rect 10115 5824 10117 5825
rect 10153 5824 10155 5825
rect 10115 5780 10116 5824
rect 10154 5780 10155 5824
rect 10115 5779 10117 5780
rect 10153 5779 10155 5780
rect 10115 5476 10117 5477
rect 10153 5476 10155 5477
rect 10115 5432 10116 5476
rect 10154 5432 10155 5476
rect 10115 5431 10117 5432
rect 10153 5431 10155 5432
rect 13116 6152 13162 6153
rect 13116 6151 13117 6152
rect 13161 6151 13162 6152
rect 13116 6114 13117 6115
rect 13161 6114 13162 6115
rect 13116 6113 13162 6114
rect 13116 5804 13162 5805
rect 13116 5803 13117 5804
rect 13161 5803 13162 5804
rect 13116 5766 13117 5767
rect 13161 5766 13162 5767
rect 13116 5765 13162 5766
rect 13116 5408 13162 5409
rect 13116 5407 13117 5408
rect 13161 5407 13162 5408
rect 13116 5370 13117 5371
rect 13161 5370 13162 5371
rect 13116 5369 13162 5370
rect 13116 5133 13162 5134
rect 13116 5132 13117 5133
rect 13161 5132 13162 5133
rect 10184 5084 13088 5085
rect 10184 5083 10185 5084
rect 13087 5083 13088 5084
rect 13116 5095 13117 5096
rect 13161 5095 13162 5096
rect 13116 5094 13162 5095
rect 10184 5054 10185 5055
rect 13087 5054 13088 5055
rect 10184 5053 13088 5054
rect 15927 3725 15929 3726
rect 15957 3725 15959 3726
rect 15927 3607 15928 3725
rect 15958 3607 15959 3725
rect 15927 3606 15929 3607
rect 15957 3606 15959 3607
<< via1 >>
rect 6452 6523 6504 6575
rect 6516 6563 6568 6575
rect 6516 6529 6522 6563
rect 6522 6529 6556 6563
rect 6556 6529 6568 6563
rect 6516 6523 6568 6529
rect 6625 6301 6805 6417
rect 13118 4859 13234 4975
rect 6776 4765 6828 4817
rect 6840 4765 6892 4817
rect 13500 3838 13680 3954
rect 13500 3774 13616 3838
rect 6452 3343 6568 3459
rect 13882 3375 13934 3427
rect 13818 3311 13870 3363
rect 13882 3311 13934 3363
rect 13112 3095 13164 3147
rect 13112 3031 13164 3083
rect 13216 3045 13268 3097
rect 13280 3045 13332 3097
rect 13286 2955 13338 3007
rect 13286 2891 13338 2943
rect 12962 2736 13078 2852
rect 13372 2580 13488 2696
rect 17108 2569 17160 2621
rect 17108 2505 17160 2557
rect 10697 2234 10877 2350
rect 17108 1754 17160 1806
rect 17108 1690 17160 1742
rect 13286 1565 13338 1617
rect 10841 1495 10893 1547
rect 10905 1495 10957 1547
rect 13286 1501 13338 1553
rect 13112 1392 13118 1426
rect 13118 1392 13152 1426
rect 13152 1392 13164 1426
rect 13112 1374 13164 1392
rect 10691 1142 10807 1322
rect 13112 1310 13164 1362
rect 13448 1089 13500 1141
rect 13448 945 13500 997
rect 13448 657 13500 709
rect 13448 513 13500 565
rect 15111 559 15163 611
rect 15111 495 15163 547
rect 17108 615 17160 667
rect 17108 551 17160 603
rect 18107 236 18159 288
rect 18171 236 18223 288
rect 13824 156 13876 208
rect 13917 156 13969 208
rect 14010 156 14062 208
rect 15117 155 15169 207
rect 13824 124 13876 144
rect 13917 124 13969 144
rect 14010 124 14062 144
rect 15117 124 15169 143
rect 17214 124 17330 208
rect 13824 92 13825 124
rect 13825 92 13859 124
rect 13859 92 13876 124
rect 13917 92 13931 124
rect 13931 92 13969 124
rect 14010 92 14041 124
rect 14041 92 14062 124
rect 15117 91 15134 124
rect 15134 91 15168 124
rect 15168 91 15169 124
rect 17214 92 17251 124
rect 17251 92 17285 124
rect 17285 92 17324 124
rect 17324 92 17330 124
<< metal2 >>
rect 6843 6575 6971 7111
rect 6446 6523 6452 6575
rect 6504 6523 6516 6575
rect 6568 6523 6574 6575
rect 6446 3459 6574 6523
rect 6602 6301 6625 6417
rect 6805 6301 6811 6417
rect 6602 4859 6811 6301
tri 6818 4817 6843 4842 se
rect 6843 4817 6898 6575
tri 6898 6550 6923 6575 nw
rect 6770 4765 6776 4817
rect 6828 4765 6840 4817
rect 6892 4765 6898 4817
rect 6926 4463 7118 5289
rect 6446 3343 6452 3459
rect 6568 3343 6574 3459
rect 12892 2852 13084 5776
rect 13112 4859 13118 4975
rect 13234 4859 13240 4975
rect 13112 4344 13240 4859
tri 13112 4216 13240 4344 ne
tri 13240 4326 13312 4398 sw
rect 13240 4216 13312 4326
tri 13240 4144 13312 4216 ne
tri 13312 4144 13494 4326 sw
tri 13312 4090 13366 4144 ne
rect 13366 3954 13494 4144
tri 13494 3954 13684 4144 sw
rect 13366 3774 13500 3954
rect 13680 3838 13686 3954
rect 13616 3774 13622 3838
tri 13622 3774 13686 3838 nw
rect 12892 2736 12962 2852
rect 13078 2736 13084 2852
rect 10691 2234 10697 2350
rect 10877 2234 10883 2350
rect 10691 1322 10807 2234
tri 10807 2158 10883 2234 nw
rect 12892 2086 13084 2736
rect 13112 3147 13164 3153
rect 13112 3083 13164 3095
rect 10691 1136 10807 1142
rect 10835 1495 10841 1547
rect 10893 1495 10905 1547
rect 10957 1495 10963 1547
rect 10835 -99 10887 1495
tri 10887 1470 10912 1495 nw
rect 13112 1426 13164 3031
rect 13112 1362 13164 1374
rect 13112 1304 13164 1310
rect 13200 3045 13216 3097
rect 13268 3045 13280 3097
rect 13332 3045 13338 3097
tri 13158 288 13200 330 se
rect 13200 308 13252 3045
tri 13252 3020 13277 3045 nw
rect 13286 3007 13338 3013
rect 13286 2943 13338 2955
rect 13286 1617 13338 2891
rect 13366 2696 13494 3774
tri 13494 3646 13622 3774 nw
tri 13841 3427 13905 3491 se
rect 13905 3427 14196 3491
tri 13789 3375 13841 3427 se
rect 13841 3375 13882 3427
rect 13934 3375 14196 3427
tri 13777 3363 13789 3375 se
rect 13789 3363 14196 3375
tri 13725 3311 13777 3363 se
rect 13777 3311 13818 3363
rect 13870 3311 13882 3363
rect 13934 3311 14196 3363
rect 13366 2580 13372 2696
rect 13488 2580 13494 2696
tri 13534 3120 13725 3311 se
rect 13725 3120 13924 3311
tri 13924 3120 14115 3311 nw
rect 13286 1553 13338 1565
rect 13286 1495 13338 1501
rect 13442 1089 13448 1141
rect 13500 1089 13506 1141
rect 13442 997 13506 1089
rect 13442 945 13448 997
rect 13500 945 13506 997
rect 13442 657 13448 709
rect 13500 657 13506 709
rect 13442 565 13506 657
rect 13442 513 13448 565
rect 13500 513 13506 565
rect 13534 462 13790 3120
tri 13790 2986 13924 3120 nw
rect 13200 288 13232 308
tri 13232 288 13252 308 nw
tri 13126 256 13158 288 se
rect 13158 256 13200 288
tri 13200 256 13232 288 nw
tri 13106 236 13126 256 se
rect 13126 236 13180 256
tri 13180 236 13200 256 nw
tri 13078 208 13106 236 se
rect 13106 208 13152 236
tri 13152 208 13180 236 nw
rect 13818 208 14074 2771
rect 15111 611 15163 617
rect 15111 547 15163 559
rect 14859 412 15052 456
tri 13052 182 13078 208 se
rect 13078 182 13126 208
tri 13126 182 13152 208 nw
tri 13026 156 13052 182 se
rect 13052 156 13100 182
tri 13100 156 13126 182 nw
rect 13818 156 13824 208
rect 13876 156 13917 208
rect 13969 156 14010 208
rect 14062 156 14074 208
tri 13025 155 13026 156 se
rect 13026 155 13099 156
tri 13099 155 13100 156 nw
tri 13014 144 13025 155 se
rect 13025 144 13088 155
tri 13088 144 13099 155 nw
rect 13818 144 14074 156
tri 12988 118 13014 144 se
rect 13014 118 13062 144
tri 13062 118 13088 144 nw
rect 12988 90 13040 118
tri 13040 96 13062 118 nw
rect 13818 92 13824 144
rect 13876 92 13917 144
rect 13969 92 14010 144
rect 14062 92 14074 144
rect 15111 208 15163 495
rect 15793 469 16113 4030
rect 17108 2621 17160 2627
rect 17108 2557 17160 2569
rect 17108 2499 17160 2505
rect 17108 1806 17160 1812
rect 17108 1742 17160 1754
rect 17108 1684 17160 1690
rect 17473 1086 17793 3504
rect 17899 3261 18219 4962
tri 17473 827 17732 1086 ne
rect 17108 667 17160 673
rect 17108 603 17160 615
rect 17108 545 17160 551
rect 17732 515 17793 1086
rect 18101 236 18107 288
rect 18159 236 18171 288
rect 18223 236 18229 288
tri 15163 208 15174 219 sw
rect 15111 207 15174 208
tri 15174 207 15175 208 sw
rect 15111 155 15117 207
rect 15169 155 15175 207
rect 15111 143 15175 155
rect 15111 91 15117 143
rect 15169 91 15175 143
rect 17208 92 17214 208
rect 17330 92 17336 208
use L1M1_CDNS_5246887918525  L1M1_CDNS_5246887918525_0
timestamp 1704896540
transform 1 0 16924 0 1 3612
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_0
timestamp 1704896540
transform 0 -1 6556 1 0 6457
box 0 0 1 1
use L1M1_CDNS_5246887918527  L1M1_CDNS_5246887918527_1
timestamp 1704896540
transform 0 -1 5826 1 0 6457
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_0
timestamp 1704896540
transform 1 0 16199 0 1 3686
box 0 0 1 1
use L1M1_CDNS_52468879185501  L1M1_CDNS_52468879185501_1
timestamp 1704896540
transform 1 0 16551 0 1 3686
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_0
timestamp 1704896540
transform 0 1 17108 -1 0 2627
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_1
timestamp 1704896540
transform 0 1 17108 -1 0 1812
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_2
timestamp 1704896540
transform 0 1 17108 -1 0 673
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_3
timestamp 1704896540
transform 0 1 13286 -1 0 3013
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_4
timestamp 1704896540
transform 0 1 13112 -1 0 1432
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_5
timestamp 1704896540
transform 0 1 13112 -1 0 3153
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_6
timestamp 1704896540
transform 0 1 13286 -1 0 1623
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_7
timestamp 1704896540
transform 0 1 15111 -1 0 617
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_8
timestamp 1704896540
transform -1 0 18229 0 1 236
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_9
timestamp 1704896540
transform -1 0 13338 0 -1 3097
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_10
timestamp 1704896540
transform -1 0 6574 0 -1 6575
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_11
timestamp 1704896540
transform 1 0 6770 0 1 4765
box 0 0 1 1
use M1M2_CDNS_5246887918577  M1M2_CDNS_5246887918577_12
timestamp 1704896540
transform 1 0 10835 0 1 1495
box 0 0 1 1
use M1M2_CDNS_52468879185197  M1M2_CDNS_52468879185197_0
timestamp 1704896540
transform 1 0 11580 0 -1 2747
box 0 0 256 116
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_0
timestamp 1704896540
transform -1 0 10883 0 -1 2350
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_1
timestamp 1704896540
transform 0 -1 10807 1 0 1136
box 0 0 1 1
use M1M2_CDNS_52468879185198  M1M2_CDNS_52468879185198_2
timestamp 1704896540
transform 1 0 6619 0 1 6301
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_0
timestamp 1704896540
transform -1 0 17336 0 1 92
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_1
timestamp 1704896540
transform -1 0 6574 0 1 3343
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_2
timestamp 1704896540
transform -1 0 13084 0 1 2736
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_3
timestamp 1704896540
transform 1 0 13366 0 -1 2696
box 0 0 1 1
use M1M2_CDNS_52468879185199  M1M2_CDNS_52468879185199_4
timestamp 1704896540
transform 1 0 13112 0 -1 4975
box 0 0 1 1
use M1M2_CDNS_52468879185200  M1M2_CDNS_52468879185200_0
timestamp 1704896540
transform 1 0 13494 0 1 3774
box 0 0 1 1
use M1M2_CDNS_52468879185201  M1M2_CDNS_52468879185201_0
timestamp 1704896540
transform 1 0 15793 0 -1 2940
box 0 0 320 116
use M1M2_CDNS_52468879185207  M1M2_CDNS_52468879185207_0
timestamp 1704896540
transform 1 0 12892 0 -1 5956
box 0 0 192 692
use M1M2_CDNS_52468879185207  M1M2_CDNS_52468879185207_1
timestamp 1704896540
transform 1 0 6926 0 1 5289
box 0 0 192 692
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_0
timestamp 1704896540
transform -1 0 13940 0 1 3311
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_1
timestamp 1704896540
transform -1 0 15175 0 1 91
box 0 0 1 1
use M1M2_CDNS_52468879185369  M1M2_CDNS_52468879185369_2
timestamp 1704896540
transform 1 0 13622 0 -1 3954
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_0
timestamp 1704896540
transform -1 0 13876 0 1 3311
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_1
timestamp 1704896540
transform 1 0 13442 0 1 1089
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_2
timestamp 1704896540
transform 1 0 13442 0 1 945
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_3
timestamp 1704896540
transform 1 0 13442 0 1 657
box 0 0 1 1
use M1M2_CDNS_52468879185970  M1M2_CDNS_52468879185970_4
timestamp 1704896540
transform 1 0 13442 0 1 513
box 0 0 1 1
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_0
timestamp 1704896540
transform 0 -1 13072 1 0 2094
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_1
timestamp 1704896540
transform 1 0 6926 0 -1 4463
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_2
timestamp 1704896540
transform 1 0 12892 0 -1 4463
box 0 0 192 180
use M1M2_CDNS_52468879185975  M1M2_CDNS_52468879185975_3
timestamp 1704896540
transform 1 0 6619 0 1 4859
box 0 0 192 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_0
timestamp 1704896540
transform 1 0 17473 0 1 3307
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_1
timestamp 1704896540
transform 1 0 17899 0 1 3307
box 0 0 320 180
use M1M2_CDNS_524688791851077  M1M2_CDNS_524688791851077_2
timestamp 1704896540
transform 1 0 17899 0 1 4769
box 0 0 320 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_0
timestamp 1704896540
transform -1 0 14196 0 1 3311
box 0 0 256 180
use M1M2_CDNS_524688791851081  M1M2_CDNS_524688791851081_1
timestamp 1704896540
transform 1 0 11580 0 -1 2050
box 0 0 256 180
use M1M2_CDNS_524688791851185  M1M2_CDNS_524688791851185_0
timestamp 1704896540
transform 1 0 15793 0 -1 4012
box 0 0 320 244
use M1M2_CDNS_524688791851458  M1M2_CDNS_524688791851458_0
timestamp 1704896540
transform 1 0 15825 0 -1 2796
box 0 0 192 2292
use M1M2_CDNS_524688791851459  M1M2_CDNS_524688791851459_0
timestamp 1704896540
transform 0 1 17732 -1 0 2627
box 0 0 2112 52
use pfet_CDNS_52468879185323  pfet_CDNS_52468879185323_0
timestamp 1704896540
transform 0 1 5874 -1 0 6622
box -119 -66 319 666
use pfet_CDNS_524688791851456  pfet_CDNS_524688791851456_0
timestamp 1704896540
transform 0 -1 13077 -1 0 5234
box -119 -66 219 3066
use pfet_CDNS_524688791851456  pfet_CDNS_524688791851456_1
timestamp 1704896540
transform 0 -1 13077 -1 0 5582
box -119 -66 219 3066
use pfet_CDNS_524688791851456  pfet_CDNS_524688791851456_2
timestamp 1704896540
transform 0 -1 13077 -1 0 5930
box -119 -66 219 3066
use pfet_CDNS_524688791851456  pfet_CDNS_524688791851456_3
timestamp 1704896540
transform 0 -1 9934 -1 0 5234
box -119 -66 219 3066
use pfet_CDNS_524688791851456  pfet_CDNS_524688791851456_4
timestamp 1704896540
transform 0 -1 9934 -1 0 5582
box -119 -66 219 3066
use pfet_CDNS_524688791851456  pfet_CDNS_524688791851456_5
timestamp 1704896540
transform 0 -1 9934 -1 0 6278
box -119 -66 219 3066
use pfet_CDNS_524688791851456  pfet_CDNS_524688791851456_6
timestamp 1704896540
transform 0 -1 9934 -1 0 5930
box -119 -66 219 3066
use pfet_CDNS_524688791851456  pfet_CDNS_524688791851456_7
timestamp 1704896540
transform 0 -1 13077 -1 0 6278
box -119 -66 219 3066
use PYL1_CDNS_52468879185444  PYL1_CDNS_52468879185444_0
timestamp 1704896540
transform 0 1 5776 1 0 6420
box 0 0 1 1
use PYL1_CDNS_524688791851460  PYL1_CDNS_524688791851460_0
timestamp 1704896540
transform 0 -1 6572 1 0 6420
box 0 0 1 1
use s8_esd_signal_5_sym_hv_local_5term  s8_esd_signal_5_sym_hv_local_5term_0
timestamp 1704896540
transform 0 -1 12948 1 0 1514
box 0 0 1591 2424
use sky130_fd_io__sio_hotswap_ctl  sky130_fd_io__sio_hotswap_ctl_0
timestamp 1704896540
transform 0 1 10691 1 0 340
box -248 -98 17453 8475
use sky130_fd_io__sio_hvsbt_inv_x1  sky130_fd_io__sio_hvsbt_inv_x1_0
timestamp 1704896540
transform -1 0 17030 0 1 3161
box -107 21 267 1369
use sky130_fd_io__sio_hvsbt_inv_x4  sky130_fd_io__sio_hvsbt_inv_x4_0
timestamp 1704896540
transform -1 0 16744 0 1 3161
box -107 21 811 1369
use sky130_fd_io__tk_em1o_b_CDNS_524688791851467  sky130_fd_io__tk_em1o_b_CDNS_524688791851467_0
timestamp 1704896540
transform 1 0 6728 0 1 5126
box 0 0 1 1
use sky130_fd_io__tk_em1o_CDNS_524688791851461  sky130_fd_io__tk_em1o_CDNS_524688791851461_0
timestamp 1704896540
transform -1 0 6652 0 -1 6417
box 0 0 1 1
use sky130_fd_io__tk_em1s_b_CDNS_524688791851463  sky130_fd_io__tk_em1s_b_CDNS_524688791851463_0
timestamp 1704896540
transform 0 -1 6892 1 0 5559
box 0 0 1 1
use sky130_fd_io__tk_em1s_b_CDNS_524688791851463  sky130_fd_io__tk_em1s_b_CDNS_524688791851463_1
timestamp 1704896540
transform 0 -1 6892 1 0 5223
box 0 0 1 1
use sky130_fd_io__tk_em1s_b_CDNS_524688791851464  sky130_fd_io__tk_em1s_b_CDNS_524688791851464_0
timestamp 1704896540
transform 0 -1 13088 1 0 5001
box 0 0 1 1
use sky130_fd_io__tk_em1s_b_CDNS_524688791851465  sky130_fd_io__tk_em1s_b_CDNS_524688791851465_0
timestamp 1704896540
transform 0 1 6920 1 0 5001
box 0 0 1 1
use sky130_fd_io__tk_em1s_b_CDNS_524688791851466  sky130_fd_io__tk_em1s_b_CDNS_524688791851466_0
timestamp 1704896540
transform -1 0 16011 0 -1 3726
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_0
timestamp 1704896540
transform -1 0 9948 0 1 6127
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_1
timestamp 1704896540
transform -1 0 9948 0 -1 5825
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_2
timestamp 1704896540
transform -1 0 9948 0 -1 5477
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_3
timestamp 1704896540
transform 1 0 10063 0 -1 5477
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_4
timestamp 1704896540
transform 1 0 10063 0 1 5779
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_52468879185341  sky130_fd_io__tk_em1s_CDNS_52468879185341_5
timestamp 1704896540
transform 1 0 10063 0 1 6127
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851462  sky130_fd_io__tk_em1s_CDNS_524688791851462_0
timestamp 1704896540
transform 0 -1 13162 -1 0 5461
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851462  sky130_fd_io__tk_em1s_CDNS_524688791851462_1
timestamp 1704896540
transform 0 -1 13162 -1 0 5857
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851462  sky130_fd_io__tk_em1s_CDNS_524688791851462_2
timestamp 1704896540
transform 0 -1 13162 -1 0 6205
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851462  sky130_fd_io__tk_em1s_CDNS_524688791851462_3
timestamp 1704896540
transform 0 1 13116 1 0 5042
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851462  sky130_fd_io__tk_em1s_CDNS_524688791851462_4
timestamp 1704896540
transform 0 1 6846 1 0 6246
box 0 0 1 1
use sky130_fd_io__tk_em1s_CDNS_524688791851462  sky130_fd_io__tk_em1s_CDNS_524688791851462_5
timestamp 1704896540
transform 0 1 6846 1 0 5989
box 0 0 1 1
<< labels >>
flabel comment s 6901 6769 6901 6769 0 FreeSans 400 90 0 0 vcc_io_soft1
flabel comment s 8450 4917 8450 4917 0 FreeSans 1400 0 0 0 pghs
flabel metal1 s 17035 3626 17035 3626 0 FreeSans 100 0 0 0 enhs_lat_h_n
flabel metal1 s 16776 4179 16776 4179 0 FreeSans 100 0 0 0 enhs_lat_h
flabel metal1 s 16368 3670 16368 3670 0 FreeSans 100 0 0 0 enhs_latbuf_h_n
flabel metal1 s 7062 4859 7254 5039 0 FreeSans 800 0 0 0 pghs_h
port 3 nsew
flabel metal1 s 5975 6523 6088 6572 0 FreeSans 400 0 0 0 padlo
port 7 nsew
flabel metal1 s 5950 6755 6373 6829 0 FreeSans 600 0 0 0 vpb_drvr
port 2 nsew
flabel metal1 s 6930 4283 7058 4463 0 FreeSans 800 0 0 0 pad
port 6 nsew
flabel metal1 s 10314 1488 10432 3315 0 FreeSans 200 0 0 0 vcc_io
port 4 nsew
flabel metal1 s 6754 5126 6778 5172 0 FreeSans 200 180 0 0 tie_hi
port 5 nsew
flabel locali s 11230 402 11578 436 0 FreeSans 200 0 0 0 vpwr_ka
port 8 nsew
flabel metal2 s 13852 92 14044 240 0 FreeSans 800 0 0 0 vgnd
port 9 nsew
flabel metal2 s 14859 412 15052 456 0 FreeSans 200 0 0 0 vcc_io
port 4 nsew
flabel metal2 s 18101 236 18229 288 0 FreeSans 200 0 0 0 od_h
port 10 nsew
flabel metal2 s 13534 466 13790 510 0 FreeSans 200 0 0 0 vgnd
port 9 nsew
flabel metal2 s 6915 7017 6915 7017 0 FreeSans 200 270 0 0 vcc_io_soft
flabel metal2 s 10835 -99 10887 -60 0 FreeSans 400 180 0 0 en_h
port 11 nsew
flabel metal2 s 12988 90 13040 112 0 FreeSans 200 0 0 0 force_h<1>
port 12 nsew
flabel nwell s 9970 5941 9994 5999 0 FreeSans 400 270 0 0 vpb_drvr
port 2 nsew
<< properties >>
string GDS_END 89236944
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 88816094
string path 345.450 3.750 351.700 3.750 
<< end >>
